//Generate the verilog at 2025-10-03T10:42:24
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00_ ;
wire _01_ ;
wire _02_ ;
wire _03_ ;
wire _04_ ;
wire _05_ ;
wire _06_ ;
wire EXU_ready_IDU ;
wire EXU_valid_LSU ;
wire EX_LS_CSRegWrite ;
wire EX_LS_RegWrite ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire IFU_valid_IDU ;
wire LSU_arready_set ;
wire LSU_awready_set ;
wire LSU_ready_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire arready_IFU ;
wire arready_LSU ;
wire arready_clint ;
wire arvalid_IFU ;
wire arvalid_LSU ;
wire arvalid_clint ;
wire awready_LSU ;
wire awvalid_LSU ;
wire bready_LSU ;
wire bvalid_LSU ;
wire check_assert ;
wire check_quest ;
wire fc_disenable ;
wire loaduse_clear ;
wire previous_load_done ;
wire rlast_IFU ;
wire rlast_LSU ;
wire rlast_clint ;
wire rmem_quest_IFU ;
wire rmem_quest_LSU ;
wire rready_IFU ;
wire rready_LSU ;
wire rready_clint ;
wire rvalid_IFU ;
wire rvalid_LSU ;
wire rvalid_clint ;
wire stall_quest_fencei ;
wire stall_quest_loaduse ;
wire wlast_LSU ;
wire wready_LSU ;
wire wvalid_LSU ;
wire \myclint/_0000_ ;
wire \myclint/_0001_ ;
wire \myclint/_0002_ ;
wire \myclint/_0003_ ;
wire \myclint/_0004_ ;
wire \myclint/_0005_ ;
wire \myclint/_0006_ ;
wire \myclint/_0007_ ;
wire \myclint/_0008_ ;
wire \myclint/_0009_ ;
wire \myclint/_0010_ ;
wire \myclint/_0011_ ;
wire \myclint/_0012_ ;
wire \myclint/_0013_ ;
wire \myclint/_0014_ ;
wire \myclint/_0015_ ;
wire \myclint/_0016_ ;
wire \myclint/_0017_ ;
wire \myclint/_0018_ ;
wire \myclint/_0019_ ;
wire \myclint/_0020_ ;
wire \myclint/_0021_ ;
wire \myclint/_0022_ ;
wire \myclint/_0023_ ;
wire \myclint/_0024_ ;
wire \myclint/_0025_ ;
wire \myclint/_0026_ ;
wire \myclint/_0027_ ;
wire \myclint/_0028_ ;
wire \myclint/_0029_ ;
wire \myclint/_0030_ ;
wire \myclint/_0031_ ;
wire \myclint/_0032_ ;
wire \myclint/_0033_ ;
wire \myclint/_0034_ ;
wire \myclint/_0035_ ;
wire \myclint/_0036_ ;
wire \myclint/_0037_ ;
wire \myclint/_0038_ ;
wire \myclint/_0039_ ;
wire \myclint/_0040_ ;
wire \myclint/_0041_ ;
wire \myclint/_0042_ ;
wire \myclint/_0043_ ;
wire \myclint/_0044_ ;
wire \myclint/_0045_ ;
wire \myclint/_0046_ ;
wire \myclint/_0047_ ;
wire \myclint/_0048_ ;
wire \myclint/_0049_ ;
wire \myclint/_0050_ ;
wire \myclint/_0051_ ;
wire \myclint/_0052_ ;
wire \myclint/_0053_ ;
wire \myclint/_0054_ ;
wire \myclint/_0055_ ;
wire \myclint/_0056_ ;
wire \myclint/_0057_ ;
wire \myclint/_0058_ ;
wire \myclint/_0059_ ;
wire \myclint/_0060_ ;
wire \myclint/_0061_ ;
wire \myclint/_0062_ ;
wire \myclint/_0063_ ;
wire \myclint/_0064_ ;
wire \myclint/_0065_ ;
wire \myclint/_0066_ ;
wire \myclint/_0067_ ;
wire \myclint/_0068_ ;
wire \myclint/_0069_ ;
wire \myclint/_0070_ ;
wire \myclint/_0071_ ;
wire \myclint/_0072_ ;
wire \myclint/_0073_ ;
wire \myclint/_0074_ ;
wire \myclint/_0075_ ;
wire \myclint/_0076_ ;
wire \myclint/_0077_ ;
wire \myclint/_0078_ ;
wire \myclint/_0079_ ;
wire \myclint/_0080_ ;
wire \myclint/_0081_ ;
wire \myclint/_0082_ ;
wire \myclint/_0083_ ;
wire \myclint/_0084_ ;
wire \myclint/_0085_ ;
wire \myclint/_0086_ ;
wire \myclint/_0087_ ;
wire \myclint/_0088_ ;
wire \myclint/_0089_ ;
wire \myclint/_0090_ ;
wire \myclint/_0091_ ;
wire \myclint/_0092_ ;
wire \myclint/_0093_ ;
wire \myclint/_0094_ ;
wire \myclint/_0095_ ;
wire \myclint/_0096_ ;
wire \myclint/_0097_ ;
wire \myclint/_0098_ ;
wire \myclint/_0099_ ;
wire \myclint/_0100_ ;
wire \myclint/_0101_ ;
wire \myclint/_0102_ ;
wire \myclint/_0103_ ;
wire \myclint/_0104_ ;
wire \myclint/_0105_ ;
wire \myclint/_0106_ ;
wire \myclint/_0107_ ;
wire \myclint/_0108_ ;
wire \myclint/_0109_ ;
wire \myclint/_0110_ ;
wire \myclint/_0111_ ;
wire \myclint/_0112_ ;
wire \myclint/_0113_ ;
wire \myclint/_0114_ ;
wire \myclint/_0115_ ;
wire \myclint/_0116_ ;
wire \myclint/_0117_ ;
wire \myclint/_0118_ ;
wire \myclint/_0119_ ;
wire \myclint/_0120_ ;
wire \myclint/_0121_ ;
wire \myclint/_0122_ ;
wire \myclint/_0123_ ;
wire \myclint/_0124_ ;
wire \myclint/_0125_ ;
wire \myclint/_0126_ ;
wire \myclint/_0127_ ;
wire \myclint/_0128_ ;
wire \myclint/_0129_ ;
wire \myclint/_0130_ ;
wire \myclint/_0131_ ;
wire \myclint/_0132_ ;
wire \myclint/_0133_ ;
wire \myclint/_0134_ ;
wire \myclint/_0135_ ;
wire \myclint/_0136_ ;
wire \myclint/_0137_ ;
wire \myclint/_0138_ ;
wire \myclint/_0139_ ;
wire \myclint/_0140_ ;
wire \myclint/_0141_ ;
wire \myclint/_0142_ ;
wire \myclint/_0143_ ;
wire \myclint/_0144_ ;
wire \myclint/_0145_ ;
wire \myclint/_0146_ ;
wire \myclint/_0147_ ;
wire \myclint/_0148_ ;
wire \myclint/_0149_ ;
wire \myclint/_0150_ ;
wire \myclint/_0151_ ;
wire \myclint/_0152_ ;
wire \myclint/_0153_ ;
wire \myclint/_0154_ ;
wire \myclint/_0155_ ;
wire \myclint/_0156_ ;
wire \myclint/_0157_ ;
wire \myclint/_0158_ ;
wire \myclint/_0159_ ;
wire \myclint/_0160_ ;
wire \myclint/_0161_ ;
wire \myclint/_0162_ ;
wire \myclint/_0163_ ;
wire \myclint/_0164_ ;
wire \myclint/_0165_ ;
wire \myclint/_0166_ ;
wire \myclint/_0167_ ;
wire \myclint/_0168_ ;
wire \myclint/_0169_ ;
wire \myclint/_0170_ ;
wire \myclint/_0171_ ;
wire \myclint/_0172_ ;
wire \myclint/_0173_ ;
wire \myclint/_0174_ ;
wire \myclint/_0175_ ;
wire \myclint/_0176_ ;
wire \myclint/_0177_ ;
wire \myclint/_0178_ ;
wire \myclint/_0179_ ;
wire \myclint/_0180_ ;
wire \myclint/_0181_ ;
wire \myclint/_0182_ ;
wire \myclint/_0183_ ;
wire \myclint/_0184_ ;
wire \myclint/_0185_ ;
wire \myclint/_0186_ ;
wire \myclint/_0187_ ;
wire \myclint/_0188_ ;
wire \myclint/_0189_ ;
wire \myclint/_0190_ ;
wire \myclint/_0191_ ;
wire \myclint/_0192_ ;
wire \myclint/_0193_ ;
wire \myclint/_0194_ ;
wire \myclint/_0195_ ;
wire \myclint/_0196_ ;
wire \myclint/_0197_ ;
wire \myclint/_0198_ ;
wire \myclint/_0199_ ;
wire \myclint/_0200_ ;
wire \myclint/_0201_ ;
wire \myclint/_0202_ ;
wire \myclint/_0203_ ;
wire \myclint/_0204_ ;
wire \myclint/_0205_ ;
wire \myclint/_0206_ ;
wire \myclint/_0207_ ;
wire \myclint/_0208_ ;
wire \myclint/_0209_ ;
wire \myclint/_0210_ ;
wire \myclint/_0211_ ;
wire \myclint/_0212_ ;
wire \myclint/_0213_ ;
wire \myclint/_0214_ ;
wire \myclint/_0215_ ;
wire \myclint/_0216_ ;
wire \myclint/_0217_ ;
wire \myclint/_0218_ ;
wire \myclint/_0219_ ;
wire \myclint/_0220_ ;
wire \myclint/_0221_ ;
wire \myclint/_0222_ ;
wire \myclint/_0223_ ;
wire \myclint/_0224_ ;
wire \myclint/_0225_ ;
wire \myclint/_0226_ ;
wire \myclint/_0227_ ;
wire \myclint/_0228_ ;
wire \myclint/_0229_ ;
wire \myclint/_0230_ ;
wire \myclint/_0231_ ;
wire \myclint/_0232_ ;
wire \myclint/_0233_ ;
wire \myclint/_0234_ ;
wire \myclint/_0235_ ;
wire \myclint/_0236_ ;
wire \myclint/_0237_ ;
wire \myclint/_0238_ ;
wire \myclint/_0239_ ;
wire \myclint/_0240_ ;
wire \myclint/_0241_ ;
wire \myclint/_0242_ ;
wire \myclint/_0243_ ;
wire \myclint/_0244_ ;
wire \myclint/_0245_ ;
wire \myclint/_0246_ ;
wire \myclint/_0247_ ;
wire \myclint/_0248_ ;
wire \myclint/_0249_ ;
wire \myclint/_0250_ ;
wire \myclint/_0251_ ;
wire \myclint/_0252_ ;
wire \myclint/_0253_ ;
wire \myclint/_0254_ ;
wire \myclint/_0255_ ;
wire \myclint/_0256_ ;
wire \myclint/_0257_ ;
wire \myclint/_0258_ ;
wire \myclint/_0259_ ;
wire \myclint/_0260_ ;
wire \myclint/_0261_ ;
wire \myclint/_0262_ ;
wire \myclint/_0263_ ;
wire \myclint/_0264_ ;
wire \myclint/_0265_ ;
wire \myclint/_0266_ ;
wire \myclint/_0267_ ;
wire \myclint/_0268_ ;
wire \myclint/_0269_ ;
wire \myclint/_0270_ ;
wire \myclint/_0271_ ;
wire \myclint/_0272_ ;
wire \myclint/_0273_ ;
wire \myclint/_0274_ ;
wire \myclint/_0275_ ;
wire \myclint/_0276_ ;
wire \myclint/_0277_ ;
wire \myclint/_0278_ ;
wire \myclint/_0279_ ;
wire \myclint/_0280_ ;
wire \myclint/_0281_ ;
wire \myclint/_0282_ ;
wire \myclint/_0283_ ;
wire \myclint/_0284_ ;
wire \myclint/_0285_ ;
wire \myclint/_0286_ ;
wire \myclint/_0287_ ;
wire \myclint/_0288_ ;
wire \myclint/_0289_ ;
wire \myclint/_0290_ ;
wire \myclint/_0291_ ;
wire \myclint/_0292_ ;
wire \myclint/_0293_ ;
wire \myclint/_0294_ ;
wire \myclint/_0295_ ;
wire \myclint/_0296_ ;
wire \myclint/_0297_ ;
wire \myclint/_0298_ ;
wire \myclint/_0299_ ;
wire \myclint/_0300_ ;
wire \myclint/_0301_ ;
wire \myclint/_0302_ ;
wire \myclint/_0303_ ;
wire \myclint/_0304_ ;
wire \myclint/_0305_ ;
wire \myclint/_0306_ ;
wire \myclint/_0307_ ;
wire \myclint/_0308_ ;
wire \myclint/_0309_ ;
wire \myclint/_0310_ ;
wire \myclint/_0311_ ;
wire \myclint/_0312_ ;
wire \myclint/_0313_ ;
wire \myclint/_0314_ ;
wire \myclint/_0315_ ;
wire \myclint/_0316_ ;
wire \myclint/_0317_ ;
wire \myclint/_0318_ ;
wire \myclint/_0319_ ;
wire \myclint/_0320_ ;
wire \myclint/_0321_ ;
wire \myclint/_0322_ ;
wire \myclint/_0323_ ;
wire \myclint/_0324_ ;
wire \myclint/_0325_ ;
wire \myclint/_0326_ ;
wire \myclint/_0327_ ;
wire \myclint/_0328_ ;
wire \myclint/_0329_ ;
wire \myclint/_0330_ ;
wire \myclint/_0331_ ;
wire \myclint/_0332_ ;
wire \myclint/_0333_ ;
wire \myclint/_0334_ ;
wire \myclint/_0335_ ;
wire \myclint/_0336_ ;
wire \myclint/_0337_ ;
wire \myclint/_0338_ ;
wire \myclint/_0339_ ;
wire \myclint/_0340_ ;
wire \myclint/_0341_ ;
wire \myclint/_0342_ ;
wire \myclint/_0343_ ;
wire \myclint/_0344_ ;
wire \myclint/_0345_ ;
wire \myclint/_0346_ ;
wire \myclint/_0347_ ;
wire \myclint/_0348_ ;
wire \myclint/_0349_ ;
wire \myclint/_0350_ ;
wire \myclint/_0351_ ;
wire \myclint/_0352_ ;
wire \myclint/_0353_ ;
wire \myclint/_0354_ ;
wire \myclint/_0355_ ;
wire \myclint/_0356_ ;
wire \myclint/_0357_ ;
wire \myclint/_0358_ ;
wire \myclint/_0359_ ;
wire \myclint/_0360_ ;
wire \myclint/_0361_ ;
wire \myclint/_0362_ ;
wire \myclint/_0363_ ;
wire \myclint/_0364_ ;
wire \myclint/_0365_ ;
wire \myclint/_0366_ ;
wire \myclint/_0367_ ;
wire \myclint/_0368_ ;
wire \myclint/_0369_ ;
wire \myclint/_0370_ ;
wire \myclint/_0371_ ;
wire \myclint/_0372_ ;
wire \myclint/_0373_ ;
wire \myclint/_0374_ ;
wire \myclint/_0375_ ;
wire \myclint/_0376_ ;
wire \myclint/_0377_ ;
wire \myclint/_0378_ ;
wire \myclint/_0379_ ;
wire \myclint/_0380_ ;
wire \myclint/_0381_ ;
wire \myclint/_0382_ ;
wire \myclint/_0383_ ;
wire \myclint/_0384_ ;
wire \myclint/_0385_ ;
wire \myclint/_0386_ ;
wire \myclint/_0387_ ;
wire \myclint/_0388_ ;
wire \myclint/_0389_ ;
wire \myclint/_0390_ ;
wire \myclint/_0391_ ;
wire \myclint/_0392_ ;
wire \myclint/_0393_ ;
wire \myclint/_0394_ ;
wire \myclint/_0395_ ;
wire \myclint/_0396_ ;
wire \myclint/_0397_ ;
wire \myclint/_0398_ ;
wire \myclint/_0399_ ;
wire \myclint/_0400_ ;
wire \myclint/_0401_ ;
wire \myclint/_0402_ ;
wire \myclint/_0403_ ;
wire \myclint/_0404_ ;
wire \myclint/_0405_ ;
wire \myclint/_0406_ ;
wire \myclint/_0407_ ;
wire \myclint/_0408_ ;
wire \myclint/_0409_ ;
wire \myclint/_0410_ ;
wire \myclint/_0411_ ;
wire \myclint/_0412_ ;
wire \myclint/_0413_ ;
wire \myclint/_0414_ ;
wire \myclint/_0415_ ;
wire \myclint/_0416_ ;
wire \myclint/_0417_ ;
wire \myclint/_0418_ ;
wire \myclint/_0419_ ;
wire \myclint/_0420_ ;
wire \myclint/_0421_ ;
wire \myclint/_0422_ ;
wire \myclint/_0423_ ;
wire \myclint/_0424_ ;
wire \myclint/_0425_ ;
wire \myclint/_0426_ ;
wire \myclint/_0427_ ;
wire \myclint/_0428_ ;
wire \myclint/_0429_ ;
wire \myclint/_0430_ ;
wire \myclint/_0431_ ;
wire \myclint/_0432_ ;
wire \myclint/_0433_ ;
wire \myclint/_0434_ ;
wire \myclint/_0435_ ;
wire \myclint/_0436_ ;
wire \myclint/_0437_ ;
wire \myclint/_0438_ ;
wire \myclint/_0439_ ;
wire \myclint/_0440_ ;
wire \myclint/_0441_ ;
wire \myclint/_0442_ ;
wire \myclint/_0443_ ;
wire \myclint/_0444_ ;
wire \myclint/_0445_ ;
wire \myclint/_0446_ ;
wire \myclint/_0447_ ;
wire \myclint/_0448_ ;
wire \myclint/_0449_ ;
wire \myclint/_0450_ ;
wire \myclint/_0451_ ;
wire \myclint/_0452_ ;
wire \myclint/_0453_ ;
wire \myclint/_0454_ ;
wire \myclint/_0455_ ;
wire \myclint/_0456_ ;
wire \myclint/_0457_ ;
wire \myclint/_0458_ ;
wire \myclint/_0459_ ;
wire \myclint/_0460_ ;
wire \myclint/_0461_ ;
wire \myclint/_0462_ ;
wire \myclint/_0463_ ;
wire \myclint/_0464_ ;
wire \myclint/_0465_ ;
wire \myclint/_0466_ ;
wire \myclint/_0467_ ;
wire \myclint/_0468_ ;
wire \myclint/_0469_ ;
wire \myclint/_0470_ ;
wire \myclint/_0471_ ;
wire \myclint/_0472_ ;
wire \myclint/_0473_ ;
wire \myclint/_0474_ ;
wire \myclint/_0475_ ;
wire \myclint/_0476_ ;
wire \myclint/_0477_ ;
wire \myclint/_0478_ ;
wire \myclint/_0479_ ;
wire \myclint/_0480_ ;
wire \myclint/_0481_ ;
wire \myclint/_0482_ ;
wire \myclint/_0483_ ;
wire \myclint/_0484_ ;
wire \myclint/_0485_ ;
wire \myclint/_0486_ ;
wire \myclint/_0487_ ;
wire \myclint/_0488_ ;
wire \myclint/_0489_ ;
wire \myclint/_0490_ ;
wire \myclint/_0491_ ;
wire \myclint/_0492_ ;
wire \myclint/_0493_ ;
wire \myclint/_0494_ ;
wire \myclint/_0495_ ;
wire \myclint/_0496_ ;
wire \myclint/_0497_ ;
wire \myclint/_0498_ ;
wire \myclint/_0499_ ;
wire \myclint/_0500_ ;
wire \myclint/_0501_ ;
wire \myclint/_0502_ ;
wire \myclint/_0503_ ;
wire \myclint/_0504_ ;
wire \myclint/_0505_ ;
wire \myclint/_0506_ ;
wire \myclint/_0507_ ;
wire \myclint/_0508_ ;
wire \myclint/_0509_ ;
wire \myclint/_0510_ ;
wire \myclint/_0511_ ;
wire \myclint/_0512_ ;
wire \myclint/_0513_ ;
wire \myclint/_0514_ ;
wire \myclint/_0515_ ;
wire \myclint/_0516_ ;
wire \myclint/_0517_ ;
wire \myclint/_0518_ ;
wire \myclint/_0519_ ;
wire \myclint/_0520_ ;
wire \myclint/_0521_ ;
wire \myclint/_0522_ ;
wire \myclint/_0523_ ;
wire \myclint/_0524_ ;
wire \myclint/_0525_ ;
wire \mycsreg/_0000_ ;
wire \mycsreg/_0001_ ;
wire \mycsreg/_0002_ ;
wire \mycsreg/_0003_ ;
wire \mycsreg/_0004_ ;
wire \mycsreg/_0005_ ;
wire \mycsreg/_0006_ ;
wire \mycsreg/_0007_ ;
wire \mycsreg/_0008_ ;
wire \mycsreg/_0009_ ;
wire \mycsreg/_0010_ ;
wire \mycsreg/_0011_ ;
wire \mycsreg/_0012_ ;
wire \mycsreg/_0013_ ;
wire \mycsreg/_0014_ ;
wire \mycsreg/_0015_ ;
wire \mycsreg/_0016_ ;
wire \mycsreg/_0017_ ;
wire \mycsreg/_0018_ ;
wire \mycsreg/_0019_ ;
wire \mycsreg/_0020_ ;
wire \mycsreg/_0021_ ;
wire \mycsreg/_0022_ ;
wire \mycsreg/_0023_ ;
wire \mycsreg/_0024_ ;
wire \mycsreg/_0025_ ;
wire \mycsreg/_0026_ ;
wire \mycsreg/_0027_ ;
wire \mycsreg/_0028_ ;
wire \mycsreg/_0029_ ;
wire \mycsreg/_0030_ ;
wire \mycsreg/_0031_ ;
wire \mycsreg/_0032_ ;
wire \mycsreg/_0033_ ;
wire \mycsreg/_0034_ ;
wire \mycsreg/_0035_ ;
wire \mycsreg/_0036_ ;
wire \mycsreg/_0037_ ;
wire \mycsreg/_0038_ ;
wire \mycsreg/_0039_ ;
wire \mycsreg/_0040_ ;
wire \mycsreg/_0041_ ;
wire \mycsreg/_0042_ ;
wire \mycsreg/_0043_ ;
wire \mycsreg/_0044_ ;
wire \mycsreg/_0045_ ;
wire \mycsreg/_0046_ ;
wire \mycsreg/_0047_ ;
wire \mycsreg/_0048_ ;
wire \mycsreg/_0049_ ;
wire \mycsreg/_0050_ ;
wire \mycsreg/_0051_ ;
wire \mycsreg/_0052_ ;
wire \mycsreg/_0053_ ;
wire \mycsreg/_0054_ ;
wire \mycsreg/_0055_ ;
wire \mycsreg/_0056_ ;
wire \mycsreg/_0057_ ;
wire \mycsreg/_0058_ ;
wire \mycsreg/_0059_ ;
wire \mycsreg/_0060_ ;
wire \mycsreg/_0061_ ;
wire \mycsreg/_0062_ ;
wire \mycsreg/_0063_ ;
wire \mycsreg/_0064_ ;
wire \mycsreg/_0065_ ;
wire \mycsreg/_0066_ ;
wire \mycsreg/_0067_ ;
wire \mycsreg/_0068_ ;
wire \mycsreg/_0069_ ;
wire \mycsreg/_0070_ ;
wire \mycsreg/_0071_ ;
wire \mycsreg/_0072_ ;
wire \mycsreg/_0073_ ;
wire \mycsreg/_0074_ ;
wire \mycsreg/_0075_ ;
wire \mycsreg/_0076_ ;
wire \mycsreg/_0077_ ;
wire \mycsreg/_0078_ ;
wire \mycsreg/_0079_ ;
wire \mycsreg/_0080_ ;
wire \mycsreg/_0081_ ;
wire \mycsreg/_0082_ ;
wire \mycsreg/_0083_ ;
wire \mycsreg/_0084_ ;
wire \mycsreg/_0085_ ;
wire \mycsreg/_0086_ ;
wire \mycsreg/_0087_ ;
wire \mycsreg/_0088_ ;
wire \mycsreg/_0089_ ;
wire \mycsreg/_0090_ ;
wire \mycsreg/_0091_ ;
wire \mycsreg/_0092_ ;
wire \mycsreg/_0093_ ;
wire \mycsreg/_0094_ ;
wire \mycsreg/_0095_ ;
wire \mycsreg/_0096_ ;
wire \mycsreg/_0097_ ;
wire \mycsreg/_0098_ ;
wire \mycsreg/_0099_ ;
wire \mycsreg/_0100_ ;
wire \mycsreg/_0101_ ;
wire \mycsreg/_0102_ ;
wire \mycsreg/_0103_ ;
wire \mycsreg/_0104_ ;
wire \mycsreg/_0105_ ;
wire \mycsreg/_0106_ ;
wire \mycsreg/_0107_ ;
wire \mycsreg/_0108_ ;
wire \mycsreg/_0109_ ;
wire \mycsreg/_0110_ ;
wire \mycsreg/_0111_ ;
wire \mycsreg/_0112_ ;
wire \mycsreg/_0113_ ;
wire \mycsreg/_0114_ ;
wire \mycsreg/_0115_ ;
wire \mycsreg/_0116_ ;
wire \mycsreg/_0117_ ;
wire \mycsreg/_0118_ ;
wire \mycsreg/_0119_ ;
wire \mycsreg/_0120_ ;
wire \mycsreg/_0121_ ;
wire \mycsreg/_0122_ ;
wire \mycsreg/_0123_ ;
wire \mycsreg/_0124_ ;
wire \mycsreg/_0125_ ;
wire \mycsreg/_0126_ ;
wire \mycsreg/_0127_ ;
wire \mycsreg/_0128_ ;
wire \mycsreg/_0129_ ;
wire \mycsreg/_0130_ ;
wire \mycsreg/_0131_ ;
wire \mycsreg/_0132_ ;
wire \mycsreg/_0133_ ;
wire \mycsreg/_0134_ ;
wire \mycsreg/_0135_ ;
wire \mycsreg/_0136_ ;
wire \mycsreg/_0137_ ;
wire \mycsreg/_0138_ ;
wire \mycsreg/_0139_ ;
wire \mycsreg/_0140_ ;
wire \mycsreg/_0141_ ;
wire \mycsreg/_0142_ ;
wire \mycsreg/_0143_ ;
wire \mycsreg/_0144_ ;
wire \mycsreg/_0145_ ;
wire \mycsreg/_0146_ ;
wire \mycsreg/_0147_ ;
wire \mycsreg/_0148_ ;
wire \mycsreg/_0149_ ;
wire \mycsreg/_0150_ ;
wire \mycsreg/_0151_ ;
wire \mycsreg/_0152_ ;
wire \mycsreg/_0153_ ;
wire \mycsreg/_0154_ ;
wire \mycsreg/_0155_ ;
wire \mycsreg/_0156_ ;
wire \mycsreg/_0157_ ;
wire \mycsreg/_0158_ ;
wire \mycsreg/_0159_ ;
wire \mycsreg/_0160_ ;
wire \mycsreg/_0161_ ;
wire \mycsreg/_0162_ ;
wire \mycsreg/_0163_ ;
wire \mycsreg/_0164_ ;
wire \mycsreg/_0165_ ;
wire \mycsreg/_0166_ ;
wire \mycsreg/_0167_ ;
wire \mycsreg/_0168_ ;
wire \mycsreg/_0169_ ;
wire \mycsreg/_0170_ ;
wire \mycsreg/_0171_ ;
wire \mycsreg/_0172_ ;
wire \mycsreg/_0173_ ;
wire \mycsreg/_0174_ ;
wire \mycsreg/_0175_ ;
wire \mycsreg/_0176_ ;
wire \mycsreg/_0177_ ;
wire \mycsreg/_0178_ ;
wire \mycsreg/_0179_ ;
wire \mycsreg/_0180_ ;
wire \mycsreg/_0181_ ;
wire \mycsreg/_0182_ ;
wire \mycsreg/_0183_ ;
wire \mycsreg/_0184_ ;
wire \mycsreg/_0185_ ;
wire \mycsreg/_0186_ ;
wire \mycsreg/_0187_ ;
wire \mycsreg/_0188_ ;
wire \mycsreg/_0189_ ;
wire \mycsreg/_0190_ ;
wire \mycsreg/_0191_ ;
wire \mycsreg/_0192_ ;
wire \mycsreg/_0193_ ;
wire \mycsreg/_0194_ ;
wire \mycsreg/_0195_ ;
wire \mycsreg/_0196_ ;
wire \mycsreg/_0197_ ;
wire \mycsreg/_0198_ ;
wire \mycsreg/_0199_ ;
wire \mycsreg/_0200_ ;
wire \mycsreg/_0201_ ;
wire \mycsreg/_0202_ ;
wire \mycsreg/_0203_ ;
wire \mycsreg/_0204_ ;
wire \mycsreg/_0205_ ;
wire \mycsreg/_0206_ ;
wire \mycsreg/_0207_ ;
wire \mycsreg/_0208_ ;
wire \mycsreg/_0209_ ;
wire \mycsreg/_0210_ ;
wire \mycsreg/_0211_ ;
wire \mycsreg/_0212_ ;
wire \mycsreg/_0213_ ;
wire \mycsreg/_0214_ ;
wire \mycsreg/_0215_ ;
wire \mycsreg/_0216_ ;
wire \mycsreg/_0217_ ;
wire \mycsreg/_0218_ ;
wire \mycsreg/_0219_ ;
wire \mycsreg/_0220_ ;
wire \mycsreg/_0221_ ;
wire \mycsreg/_0222_ ;
wire \mycsreg/_0223_ ;
wire \mycsreg/_0224_ ;
wire \mycsreg/_0225_ ;
wire \mycsreg/_0226_ ;
wire \mycsreg/_0227_ ;
wire \mycsreg/_0228_ ;
wire \mycsreg/_0229_ ;
wire \mycsreg/_0230_ ;
wire \mycsreg/_0231_ ;
wire \mycsreg/_0232_ ;
wire \mycsreg/_0233_ ;
wire \mycsreg/_0234_ ;
wire \mycsreg/_0235_ ;
wire \mycsreg/_0236_ ;
wire \mycsreg/_0237_ ;
wire \mycsreg/_0238_ ;
wire \mycsreg/_0239_ ;
wire \mycsreg/_0240_ ;
wire \mycsreg/_0241_ ;
wire \mycsreg/_0242_ ;
wire \mycsreg/_0243_ ;
wire \mycsreg/_0244_ ;
wire \mycsreg/_0245_ ;
wire \mycsreg/_0246_ ;
wire \mycsreg/_0247_ ;
wire \mycsreg/_0248_ ;
wire \mycsreg/_0249_ ;
wire \mycsreg/_0250_ ;
wire \mycsreg/_0251_ ;
wire \mycsreg/_0252_ ;
wire \mycsreg/_0253_ ;
wire \mycsreg/_0254_ ;
wire \mycsreg/_0255_ ;
wire \mycsreg/_0256_ ;
wire \mycsreg/_0257_ ;
wire \mycsreg/_0258_ ;
wire \mycsreg/_0259_ ;
wire \mycsreg/_0260_ ;
wire \mycsreg/_0261_ ;
wire \mycsreg/_0262_ ;
wire \mycsreg/_0263_ ;
wire \mycsreg/_0264_ ;
wire \mycsreg/_0265_ ;
wire \mycsreg/_0266_ ;
wire \mycsreg/_0267_ ;
wire \mycsreg/_0268_ ;
wire \mycsreg/_0269_ ;
wire \mycsreg/_0270_ ;
wire \mycsreg/_0271_ ;
wire \mycsreg/_0272_ ;
wire \mycsreg/_0273_ ;
wire \mycsreg/_0274_ ;
wire \mycsreg/_0275_ ;
wire \mycsreg/_0276_ ;
wire \mycsreg/_0277_ ;
wire \mycsreg/_0278_ ;
wire \mycsreg/_0279_ ;
wire \mycsreg/_0280_ ;
wire \mycsreg/_0281_ ;
wire \mycsreg/_0282_ ;
wire \mycsreg/_0283_ ;
wire \mycsreg/_0284_ ;
wire \mycsreg/_0285_ ;
wire \mycsreg/_0286_ ;
wire \mycsreg/_0287_ ;
wire \mycsreg/_0288_ ;
wire \mycsreg/_0289_ ;
wire \mycsreg/_0290_ ;
wire \mycsreg/_0291_ ;
wire \mycsreg/_0292_ ;
wire \mycsreg/_0293_ ;
wire \mycsreg/_0294_ ;
wire \mycsreg/_0295_ ;
wire \mycsreg/_0296_ ;
wire \mycsreg/_0297_ ;
wire \mycsreg/_0298_ ;
wire \mycsreg/_0299_ ;
wire \mycsreg/_0300_ ;
wire \mycsreg/_0301_ ;
wire \mycsreg/_0302_ ;
wire \mycsreg/_0303_ ;
wire \mycsreg/_0304_ ;
wire \mycsreg/_0305_ ;
wire \mycsreg/_0306_ ;
wire \mycsreg/_0307_ ;
wire \mycsreg/_0308_ ;
wire \mycsreg/_0309_ ;
wire \mycsreg/_0310_ ;
wire \mycsreg/_0311_ ;
wire \mycsreg/_0312_ ;
wire \mycsreg/_0313_ ;
wire \mycsreg/_0314_ ;
wire \mycsreg/_0315_ ;
wire \mycsreg/_0316_ ;
wire \mycsreg/_0317_ ;
wire \mycsreg/_0318_ ;
wire \mycsreg/_0319_ ;
wire \mycsreg/_0320_ ;
wire \mycsreg/_0321_ ;
wire \mycsreg/_0322_ ;
wire \mycsreg/_0323_ ;
wire \mycsreg/_0324_ ;
wire \mycsreg/_0325_ ;
wire \mycsreg/_0326_ ;
wire \mycsreg/_0327_ ;
wire \mycsreg/_0328_ ;
wire \mycsreg/_0329_ ;
wire \mycsreg/_0330_ ;
wire \mycsreg/_0331_ ;
wire \mycsreg/_0332_ ;
wire \mycsreg/_0333_ ;
wire \mycsreg/_0334_ ;
wire \mycsreg/_0335_ ;
wire \mycsreg/_0336_ ;
wire \mycsreg/_0337_ ;
wire \mycsreg/_0338_ ;
wire \mycsreg/_0339_ ;
wire \mycsreg/_0340_ ;
wire \mycsreg/_0341_ ;
wire \mycsreg/_0342_ ;
wire \mycsreg/_0343_ ;
wire \mycsreg/_0344_ ;
wire \mycsreg/_0345_ ;
wire \mycsreg/_0346_ ;
wire \mycsreg/_0347_ ;
wire \mycsreg/_0348_ ;
wire \mycsreg/_0349_ ;
wire \mycsreg/_0350_ ;
wire \mycsreg/_0351_ ;
wire \mycsreg/_0352_ ;
wire \mycsreg/_0353_ ;
wire \mycsreg/_0354_ ;
wire \mycsreg/_0355_ ;
wire \mycsreg/_0356_ ;
wire \mycsreg/_0357_ ;
wire \mycsreg/_0358_ ;
wire \mycsreg/_0359_ ;
wire \mycsreg/_0360_ ;
wire \mycsreg/_0361_ ;
wire \mycsreg/_0362_ ;
wire \mycsreg/_0363_ ;
wire \mycsreg/_0364_ ;
wire \mycsreg/_0365_ ;
wire \mycsreg/_0366_ ;
wire \mycsreg/_0367_ ;
wire \mycsreg/_0368_ ;
wire \mycsreg/_0369_ ;
wire \mycsreg/_0370_ ;
wire \mycsreg/_0371_ ;
wire \mycsreg/_0372_ ;
wire \mycsreg/_0373_ ;
wire \mycsreg/_0374_ ;
wire \mycsreg/_0375_ ;
wire \mycsreg/_0376_ ;
wire \mycsreg/_0377_ ;
wire \mycsreg/_0378_ ;
wire \mycsreg/_0379_ ;
wire \mycsreg/_0380_ ;
wire \mycsreg/_0381_ ;
wire \mycsreg/_0382_ ;
wire \mycsreg/_0383_ ;
wire \mycsreg/_0384_ ;
wire \mycsreg/_0385_ ;
wire \mycsreg/_0386_ ;
wire \mycsreg/_0387_ ;
wire \mycsreg/_0388_ ;
wire \mycsreg/_0389_ ;
wire \mycsreg/_0390_ ;
wire \mycsreg/_0391_ ;
wire \mycsreg/_0392_ ;
wire \mycsreg/_0393_ ;
wire \mycsreg/_0394_ ;
wire \mycsreg/_0395_ ;
wire \mycsreg/_0396_ ;
wire \mycsreg/_0397_ ;
wire \mycsreg/_0398_ ;
wire \mycsreg/_0399_ ;
wire \mycsreg/_0400_ ;
wire \mycsreg/_0401_ ;
wire \mycsreg/_0402_ ;
wire \mycsreg/_0403_ ;
wire \mycsreg/_0404_ ;
wire \mycsreg/_0405_ ;
wire \mycsreg/_0406_ ;
wire \mycsreg/_0407_ ;
wire \mycsreg/_0408_ ;
wire \mycsreg/_0409_ ;
wire \mycsreg/_0410_ ;
wire \mycsreg/_0411_ ;
wire \mycsreg/_0412_ ;
wire \mycsreg/_0413_ ;
wire \mycsreg/_0414_ ;
wire \mycsreg/_0415_ ;
wire \mycsreg/_0416_ ;
wire \mycsreg/_0417_ ;
wire \mycsreg/_0418_ ;
wire \mycsreg/_0419_ ;
wire \mycsreg/_0420_ ;
wire \mycsreg/_0421_ ;
wire \mycsreg/_0422_ ;
wire \mycsreg/_0423_ ;
wire \mycsreg/_0424_ ;
wire \mycsreg/_0425_ ;
wire \mycsreg/_0426_ ;
wire \mycsreg/_0427_ ;
wire \mycsreg/_0428_ ;
wire \mycsreg/_0429_ ;
wire \mycsreg/_0430_ ;
wire \mycsreg/_0431_ ;
wire \mycsreg/_0432_ ;
wire \mycsreg/_0433_ ;
wire \mycsreg/_0434_ ;
wire \mycsreg/_0435_ ;
wire \mycsreg/_0436_ ;
wire \mycsreg/_0437_ ;
wire \mycsreg/_0438_ ;
wire \mycsreg/_0439_ ;
wire \mycsreg/_0440_ ;
wire \mycsreg/_0441_ ;
wire \mycsreg/_0442_ ;
wire \mycsreg/_0443_ ;
wire \mycsreg/_0444_ ;
wire \mycsreg/_0445_ ;
wire \mycsreg/_0446_ ;
wire \mycsreg/_0447_ ;
wire \mycsreg/_0448_ ;
wire \mycsreg/_0449_ ;
wire \mycsreg/_0450_ ;
wire \mycsreg/_0451_ ;
wire \mycsreg/_0452_ ;
wire \mycsreg/_0453_ ;
wire \mycsreg/_0454_ ;
wire \mycsreg/_0455_ ;
wire \mycsreg/_0456_ ;
wire \mycsreg/_0457_ ;
wire \mycsreg/_0458_ ;
wire \mycsreg/_0459_ ;
wire \mycsreg/_0460_ ;
wire \mycsreg/_0461_ ;
wire \mycsreg/_0462_ ;
wire \mycsreg/_0463_ ;
wire \mycsreg/_0464_ ;
wire \mycsreg/_0465_ ;
wire \mycsreg/_0466_ ;
wire \mycsreg/_0467_ ;
wire \mycsreg/_0468_ ;
wire \mycsreg/_0469_ ;
wire \mycsreg/_0470_ ;
wire \mycsreg/_0471_ ;
wire \mycsreg/_0472_ ;
wire \mycsreg/_0473_ ;
wire \mycsreg/_0474_ ;
wire \mycsreg/_0475_ ;
wire \mycsreg/_0476_ ;
wire \mycsreg/_0477_ ;
wire \mycsreg/_0478_ ;
wire \mycsreg/_0479_ ;
wire \mycsreg/_0480_ ;
wire \mycsreg/_0481_ ;
wire \mycsreg/_0482_ ;
wire \mycsreg/_0483_ ;
wire \mycsreg/_0484_ ;
wire \mycsreg/_0485_ ;
wire \mycsreg/_0486_ ;
wire \mycsreg/_0487_ ;
wire \mycsreg/_0488_ ;
wire \mycsreg/_0489_ ;
wire \mycsreg/_0490_ ;
wire \mycsreg/_0491_ ;
wire \mycsreg/_0492_ ;
wire \mycsreg/_0493_ ;
wire \mycsreg/_0494_ ;
wire \mycsreg/_0495_ ;
wire \mycsreg/_0496_ ;
wire \mycsreg/_0497_ ;
wire \mycsreg/_0498_ ;
wire \mycsreg/_0499_ ;
wire \mycsreg/_0500_ ;
wire \mycsreg/_0501_ ;
wire \mycsreg/_0502_ ;
wire \mycsreg/_0503_ ;
wire \mycsreg/_0504_ ;
wire \mycsreg/_0505_ ;
wire \mycsreg/_0506_ ;
wire \mycsreg/_0507_ ;
wire \mycsreg/_0508_ ;
wire \mycsreg/_0509_ ;
wire \mycsreg/_0510_ ;
wire \mycsreg/_0511_ ;
wire \mycsreg/_0512_ ;
wire \mycsreg/_0513_ ;
wire \mycsreg/_0514_ ;
wire \mycsreg/_0515_ ;
wire \mycsreg/_0516_ ;
wire \mycsreg/_0517_ ;
wire \mycsreg/_0518_ ;
wire \mycsreg/_0519_ ;
wire \mycsreg/_0520_ ;
wire \mycsreg/_0521_ ;
wire \mycsreg/_0522_ ;
wire \mycsreg/_0523_ ;
wire \mycsreg/_0524_ ;
wire \mycsreg/_0525_ ;
wire \mycsreg/_0526_ ;
wire \mycsreg/_0527_ ;
wire \mycsreg/_0528_ ;
wire \mycsreg/_0529_ ;
wire \mycsreg/_0530_ ;
wire \mycsreg/_0531_ ;
wire \mycsreg/_0532_ ;
wire \mycsreg/_0533_ ;
wire \mycsreg/_0534_ ;
wire \mycsreg/_0535_ ;
wire \mycsreg/_0536_ ;
wire \mycsreg/_0537_ ;
wire \mycsreg/_0538_ ;
wire \mycsreg/_0539_ ;
wire \mycsreg/_0540_ ;
wire \mycsreg/_0541_ ;
wire \mycsreg/_0542_ ;
wire \mycsreg/_0543_ ;
wire \mycsreg/_0544_ ;
wire \mycsreg/_0545_ ;
wire \mycsreg/_0546_ ;
wire \mycsreg/_0547_ ;
wire \mycsreg/_0548_ ;
wire \mycsreg/_0549_ ;
wire \mycsreg/_0550_ ;
wire \mycsreg/_0551_ ;
wire \mycsreg/_0552_ ;
wire \mycsreg/_0553_ ;
wire \mycsreg/_0554_ ;
wire \mycsreg/_0555_ ;
wire \mycsreg/_0556_ ;
wire \mycsreg/_0557_ ;
wire \mycsreg/_0558_ ;
wire \mycsreg/_0559_ ;
wire \mycsreg/_0560_ ;
wire \mycsreg/_0561_ ;
wire \mycsreg/_0562_ ;
wire \mycsreg/_0563_ ;
wire \mycsreg/_0564_ ;
wire \mycsreg/_0565_ ;
wire \mycsreg/_0566_ ;
wire \mycsreg/_0567_ ;
wire \mycsreg/_0568_ ;
wire \mycsreg/_0569_ ;
wire \mycsreg/_0570_ ;
wire \mycsreg/_0571_ ;
wire \mycsreg/_0572_ ;
wire \mycsreg/_0573_ ;
wire \mycsreg/_0574_ ;
wire \mycsreg/_0575_ ;
wire \mycsreg/_0576_ ;
wire \mycsreg/_0577_ ;
wire \mycsreg/_0578_ ;
wire \mycsreg/_0579_ ;
wire \mycsreg/_0580_ ;
wire \mycsreg/_0581_ ;
wire \mycsreg/_0582_ ;
wire \mycsreg/_0583_ ;
wire \mycsreg/_0584_ ;
wire \mycsreg/_0585_ ;
wire \mycsreg/_0586_ ;
wire \mycsreg/_0587_ ;
wire \mycsreg/_0588_ ;
wire \mycsreg/_0589_ ;
wire \mycsreg/_0590_ ;
wire \mycsreg/_0591_ ;
wire \mycsreg/_0592_ ;
wire \mycsreg/_0593_ ;
wire \mycsreg/_0594_ ;
wire \mycsreg/_0595_ ;
wire \mycsreg/_0596_ ;
wire \mycsreg/_0597_ ;
wire \mycsreg/_0598_ ;
wire \mycsreg/_0599_ ;
wire \mycsreg/_0600_ ;
wire \mycsreg/_0601_ ;
wire \mycsreg/_0602_ ;
wire \mycsreg/_0603_ ;
wire \mycsreg/_0604_ ;
wire \mycsreg/_0605_ ;
wire \mycsreg/_0606_ ;
wire \mycsreg/_0607_ ;
wire \mycsreg/_0608_ ;
wire \mycsreg/_0609_ ;
wire \mycsreg/_0610_ ;
wire \mycsreg/_0611_ ;
wire \mycsreg/_0612_ ;
wire \mycsreg/_0613_ ;
wire \mycsreg/_0614_ ;
wire \mycsreg/_0615_ ;
wire \mycsreg/_0616_ ;
wire \mycsreg/_0617_ ;
wire \mycsreg/_0618_ ;
wire \mycsreg/_0619_ ;
wire \mycsreg/_0620_ ;
wire \mycsreg/_0621_ ;
wire \mycsreg/_0622_ ;
wire \mycsreg/_0623_ ;
wire \mycsreg/_0624_ ;
wire \mycsreg/_0625_ ;
wire \mycsreg/_0626_ ;
wire \mycsreg/_0627_ ;
wire \mycsreg/_0628_ ;
wire \mycsreg/_0629_ ;
wire \mycsreg/_0630_ ;
wire \mycsreg/_0631_ ;
wire \mycsreg/_0632_ ;
wire \mycsreg/_0633_ ;
wire \mycsreg/_0634_ ;
wire \mycsreg/_0635_ ;
wire \mycsreg/_0636_ ;
wire \mycsreg/_0637_ ;
wire \mycsreg/_0638_ ;
wire \mycsreg/_0639_ ;
wire \mycsreg/_0640_ ;
wire \mycsreg/_0641_ ;
wire \mycsreg/_0642_ ;
wire \mycsreg/_0643_ ;
wire \mycsreg/_0644_ ;
wire \mycsreg/_0645_ ;
wire \mycsreg/_0646_ ;
wire \mycsreg/_0647_ ;
wire \mycsreg/_0648_ ;
wire \mycsreg/_0649_ ;
wire \mycsreg/_0650_ ;
wire \mycsreg/_0651_ ;
wire \mycsreg/_0652_ ;
wire \mycsreg/_0653_ ;
wire \mycsreg/_0654_ ;
wire \mycsreg/_0655_ ;
wire \mycsreg/_0656_ ;
wire \mycsreg/_0657_ ;
wire \mycsreg/_0658_ ;
wire \mycsreg/_0659_ ;
wire \mycsreg/_0660_ ;
wire \mycsreg/_0661_ ;
wire \mycsreg/_0662_ ;
wire \mycsreg/_0663_ ;
wire \mycsreg/_0664_ ;
wire \mycsreg/_0665_ ;
wire \mycsreg/_0666_ ;
wire \mycsreg/_0667_ ;
wire \mycsreg/_0668_ ;
wire \mycsreg/_0669_ ;
wire \mycsreg/_0670_ ;
wire \mycsreg/_0671_ ;
wire \mycsreg/_0672_ ;
wire \mycsreg/_0673_ ;
wire \mycsreg/_0674_ ;
wire \mycsreg/_0675_ ;
wire \mycsreg/_0676_ ;
wire \mycsreg/_0677_ ;
wire \mycsreg/_0678_ ;
wire \mycsreg/_0679_ ;
wire \mycsreg/_0680_ ;
wire \mycsreg/_0681_ ;
wire \mycsreg/_0682_ ;
wire \mycsreg/_0683_ ;
wire \mycsreg/_0684_ ;
wire \mycsreg/_0685_ ;
wire \mycsreg/_0686_ ;
wire \mycsreg/_0687_ ;
wire \mycsreg/_0688_ ;
wire \mycsreg/_0689_ ;
wire \mycsreg/_0690_ ;
wire \mycsreg/_0691_ ;
wire \mycsreg/_0692_ ;
wire \mycsreg/_0693_ ;
wire \mycsreg/_0694_ ;
wire \mycsreg/_0695_ ;
wire \mycsreg/_0696_ ;
wire \mycsreg/_0697_ ;
wire \mycsreg/_0698_ ;
wire \mycsreg/_0699_ ;
wire \mycsreg/_0700_ ;
wire \mycsreg/_0701_ ;
wire \mycsreg/_0702_ ;
wire \mycsreg/_0703_ ;
wire \mycsreg/_0704_ ;
wire \mycsreg/_0705_ ;
wire \mycsreg/_0706_ ;
wire \mycsreg/_0707_ ;
wire \mycsreg/_0708_ ;
wire \mycsreg/_0709_ ;
wire \mycsreg/_0710_ ;
wire \mycsreg/_0711_ ;
wire \mycsreg/_0712_ ;
wire \mycsreg/_0713_ ;
wire \mycsreg/_0714_ ;
wire \mycsreg/_0715_ ;
wire \mycsreg/_0716_ ;
wire \mycsreg/_0717_ ;
wire \mycsreg/_0718_ ;
wire \mycsreg/_0719_ ;
wire \mycsreg/_0720_ ;
wire \mycsreg/_0721_ ;
wire \mycsreg/_0722_ ;
wire \mycsreg/_0723_ ;
wire \mycsreg/_0724_ ;
wire \mycsreg/_0725_ ;
wire \mycsreg/_0726_ ;
wire \mycsreg/_0727_ ;
wire \mycsreg/_0728_ ;
wire \mycsreg/_0729_ ;
wire \mycsreg/_0730_ ;
wire \mycsreg/_0731_ ;
wire \mycsreg/_0732_ ;
wire \mycsreg/_0733_ ;
wire \mycsreg/_0734_ ;
wire \mycsreg/_0735_ ;
wire \mycsreg/_0736_ ;
wire \mycsreg/_0737_ ;
wire \mycsreg/_0738_ ;
wire \mycsreg/_0739_ ;
wire \mycsreg/_0740_ ;
wire \mycsreg/_0741_ ;
wire \mycsreg/_0742_ ;
wire \mycsreg/_0743_ ;
wire \mycsreg/_0744_ ;
wire \mycsreg/_0745_ ;
wire \mycsreg/_0746_ ;
wire \mycsreg/_0747_ ;
wire \mycsreg/_0748_ ;
wire \mycsreg/_0749_ ;
wire \mycsreg/_0750_ ;
wire \mycsreg/_0751_ ;
wire \mycsreg/_0752_ ;
wire \mycsreg/_0753_ ;
wire \mycsreg/_0754_ ;
wire \mycsreg/_0755_ ;
wire \mycsreg/_0756_ ;
wire \mycsreg/_0757_ ;
wire \mycsreg/_0758_ ;
wire \mycsreg/_0759_ ;
wire \mycsreg/_0760_ ;
wire \mycsreg/_0761_ ;
wire \mycsreg/_0762_ ;
wire \mycsreg/_0763_ ;
wire \mycsreg/_0764_ ;
wire \mycsreg/_0765_ ;
wire \mycsreg/_0766_ ;
wire \mycsreg/_0767_ ;
wire \mycsreg/_0768_ ;
wire \mycsreg/_0769_ ;
wire \mycsreg/_0770_ ;
wire \mycsreg/_0771_ ;
wire \mycsreg/_0772_ ;
wire \mycsreg/_0773_ ;
wire \mycsreg/_0774_ ;
wire \mycsreg/_0775_ ;
wire \mycsreg/_0776_ ;
wire \mycsreg/_0777_ ;
wire \mycsreg/_0778_ ;
wire \mycsreg/_0779_ ;
wire \mycsreg/_0780_ ;
wire \mycsreg/_0781_ ;
wire \mycsreg/_0782_ ;
wire \mycsreg/_0783_ ;
wire \mycsreg/_0784_ ;
wire \mycsreg/_0785_ ;
wire \mycsreg/_0786_ ;
wire \mycsreg/_0787_ ;
wire \mycsreg/_0788_ ;
wire \mycsreg/_0789_ ;
wire \mycsreg/_0790_ ;
wire \mycsreg/_0791_ ;
wire \mycsreg/_0792_ ;
wire \mycsreg/_0793_ ;
wire \mycsreg/_0794_ ;
wire \mycsreg/_0795_ ;
wire \mycsreg/_0796_ ;
wire \mycsreg/_0797_ ;
wire \mycsreg/_0798_ ;
wire \mycsreg/_0799_ ;
wire \mycsreg/_0800_ ;
wire \mycsreg/_0801_ ;
wire \mycsreg/_0802_ ;
wire \mycsreg/_0803_ ;
wire \mycsreg/_0804_ ;
wire \mycsreg/_0805_ ;
wire \mycsreg/_0806_ ;
wire \mycsreg/_0807_ ;
wire \mycsreg/_0808_ ;
wire \mycsreg/_0809_ ;
wire \mycsreg/_0810_ ;
wire \mycsreg/_0811_ ;
wire \mycsreg/_0812_ ;
wire \mycsreg/_0813_ ;
wire \mycsreg/_0814_ ;
wire \mycsreg/_0815_ ;
wire \mycsreg/_0816_ ;
wire \mycsreg/_0817_ ;
wire \mycsreg/_0818_ ;
wire \mycsreg/_0819_ ;
wire \mycsreg/_0820_ ;
wire \mycsreg/_0821_ ;
wire \mycsreg/_0822_ ;
wire \mycsreg/_0823_ ;
wire \mycsreg/_0824_ ;
wire \mycsreg/_0825_ ;
wire \mycsreg/_0826_ ;
wire \mycsreg/_0827_ ;
wire \mycsreg/_0828_ ;
wire \mycsreg/_0829_ ;
wire \mycsreg/_0830_ ;
wire \mycsreg/_0831_ ;
wire \mycsreg/_0832_ ;
wire \mycsreg/_0833_ ;
wire \mycsreg/_0834_ ;
wire \mycsreg/_0835_ ;
wire \mycsreg/_0836_ ;
wire \mycsreg/_0837_ ;
wire \mycsreg/_0838_ ;
wire \mycsreg/_0839_ ;
wire \mycsreg/_0840_ ;
wire \mycsreg/_0841_ ;
wire \mycsreg/_0842_ ;
wire \mycsreg/_0843_ ;
wire \mycsreg/_0844_ ;
wire \mycsreg/_0845_ ;
wire \mycsreg/_0846_ ;
wire \mycsreg/_0847_ ;
wire \mycsreg/_0848_ ;
wire \mycsreg/_0849_ ;
wire \mycsreg/_0850_ ;
wire \mycsreg/_0851_ ;
wire \mycsreg/_0852_ ;
wire \mycsreg/_0853_ ;
wire \mycsreg/_0854_ ;
wire \mycsreg/_0855_ ;
wire \mycsreg/_0856_ ;
wire \mycsreg/_0857_ ;
wire \mycsreg/_0858_ ;
wire \mycsreg/_0859_ ;
wire \mycsreg/_0860_ ;
wire \mycsreg/_0861_ ;
wire \mycsreg/_0862_ ;
wire \mycsreg/_0863_ ;
wire \mycsreg/_0864_ ;
wire \mycsreg/_0865_ ;
wire \mycsreg/_0866_ ;
wire \mycsreg/_0867_ ;
wire \mycsreg/_0868_ ;
wire \mycsreg/_0869_ ;
wire \mycsreg/_0870_ ;
wire \mycsreg/_0871_ ;
wire \mycsreg/_0872_ ;
wire \mycsreg/_0873_ ;
wire \mycsreg/_0874_ ;
wire \mycsreg/_0875_ ;
wire \mycsreg/_0876_ ;
wire \mycsreg/_0877_ ;
wire \mycsreg/_0878_ ;
wire \mycsreg/_0879_ ;
wire \mycsreg/_0880_ ;
wire \mycsreg/_0881_ ;
wire \mycsreg/_0882_ ;
wire \mycsreg/_0883_ ;
wire \mycsreg/_0884_ ;
wire \mycsreg/_0885_ ;
wire \mycsreg/_0886_ ;
wire \mycsreg/_0887_ ;
wire \mycsreg/_0888_ ;
wire \mycsreg/_0889_ ;
wire \mycsreg/_0890_ ;
wire \mycsreg/_0891_ ;
wire \mycsreg/_0892_ ;
wire \mycsreg/_0893_ ;
wire \mycsreg/_0894_ ;
wire \mycsreg/_0895_ ;
wire \mycsreg/_0896_ ;
wire \mycsreg/_0897_ ;
wire \mycsreg/_0898_ ;
wire \mycsreg/_0899_ ;
wire \mycsreg/_0900_ ;
wire \mycsreg/_0901_ ;
wire \mycsreg/_0902_ ;
wire \mycsreg/_0903_ ;
wire \mycsreg/_0904_ ;
wire \mycsreg/_0905_ ;
wire \mycsreg/_0906_ ;
wire \mycsreg/_0907_ ;
wire \mycsreg/_0908_ ;
wire \mycsreg/_0909_ ;
wire \mycsreg/_0910_ ;
wire \mycsreg/_0911_ ;
wire \mycsreg/_0912_ ;
wire \mycsreg/_0913_ ;
wire \mycsreg/_0914_ ;
wire \mycsreg/_0915_ ;
wire \mycsreg/_0916_ ;
wire \mycsreg/_0917_ ;
wire \mycsreg/_0918_ ;
wire \mycsreg/_0919_ ;
wire \mycsreg/_0920_ ;
wire \mycsreg/_0921_ ;
wire \mycsreg/_0922_ ;
wire \mycsreg/_0923_ ;
wire \mycsreg/_0924_ ;
wire \mycsreg/_0925_ ;
wire \mycsreg/_0926_ ;
wire \mycsreg/_0927_ ;
wire \mycsreg/_0928_ ;
wire \mycsreg/_0929_ ;
wire \mycsreg/_0930_ ;
wire \mycsreg/_0931_ ;
wire \mycsreg/CSReg[0][0] ;
wire \mycsreg/CSReg[0][10] ;
wire \mycsreg/CSReg[0][11] ;
wire \mycsreg/CSReg[0][12] ;
wire \mycsreg/CSReg[0][13] ;
wire \mycsreg/CSReg[0][14] ;
wire \mycsreg/CSReg[0][15] ;
wire \mycsreg/CSReg[0][16] ;
wire \mycsreg/CSReg[0][17] ;
wire \mycsreg/CSReg[0][18] ;
wire \mycsreg/CSReg[0][19] ;
wire \mycsreg/CSReg[0][1] ;
wire \mycsreg/CSReg[0][20] ;
wire \mycsreg/CSReg[0][21] ;
wire \mycsreg/CSReg[0][22] ;
wire \mycsreg/CSReg[0][23] ;
wire \mycsreg/CSReg[0][24] ;
wire \mycsreg/CSReg[0][25] ;
wire \mycsreg/CSReg[0][26] ;
wire \mycsreg/CSReg[0][27] ;
wire \mycsreg/CSReg[0][28] ;
wire \mycsreg/CSReg[0][29] ;
wire \mycsreg/CSReg[0][2] ;
wire \mycsreg/CSReg[0][30] ;
wire \mycsreg/CSReg[0][31] ;
wire \mycsreg/CSReg[0][3] ;
wire \mycsreg/CSReg[0][4] ;
wire \mycsreg/CSReg[0][5] ;
wire \mycsreg/CSReg[0][6] ;
wire \mycsreg/CSReg[0][7] ;
wire \mycsreg/CSReg[0][8] ;
wire \mycsreg/CSReg[0][9] ;
wire \mycsreg/CSReg[1][0] ;
wire \mycsreg/CSReg[1][10] ;
wire \mycsreg/CSReg[1][11] ;
wire \mycsreg/CSReg[1][12] ;
wire \mycsreg/CSReg[1][13] ;
wire \mycsreg/CSReg[1][14] ;
wire \mycsreg/CSReg[1][15] ;
wire \mycsreg/CSReg[1][16] ;
wire \mycsreg/CSReg[1][17] ;
wire \mycsreg/CSReg[1][18] ;
wire \mycsreg/CSReg[1][19] ;
wire \mycsreg/CSReg[1][1] ;
wire \mycsreg/CSReg[1][20] ;
wire \mycsreg/CSReg[1][21] ;
wire \mycsreg/CSReg[1][22] ;
wire \mycsreg/CSReg[1][23] ;
wire \mycsreg/CSReg[1][24] ;
wire \mycsreg/CSReg[1][25] ;
wire \mycsreg/CSReg[1][26] ;
wire \mycsreg/CSReg[1][27] ;
wire \mycsreg/CSReg[1][28] ;
wire \mycsreg/CSReg[1][29] ;
wire \mycsreg/CSReg[1][2] ;
wire \mycsreg/CSReg[1][30] ;
wire \mycsreg/CSReg[1][31] ;
wire \mycsreg/CSReg[1][3] ;
wire \mycsreg/CSReg[1][4] ;
wire \mycsreg/CSReg[1][5] ;
wire \mycsreg/CSReg[1][6] ;
wire \mycsreg/CSReg[1][7] ;
wire \mycsreg/CSReg[1][8] ;
wire \mycsreg/CSReg[1][9] ;
wire \mycsreg/CSReg[2][0] ;
wire \mycsreg/CSReg[2][10] ;
wire \mycsreg/CSReg[2][11] ;
wire \mycsreg/CSReg[2][12] ;
wire \mycsreg/CSReg[2][13] ;
wire \mycsreg/CSReg[2][14] ;
wire \mycsreg/CSReg[2][15] ;
wire \mycsreg/CSReg[2][16] ;
wire \mycsreg/CSReg[2][17] ;
wire \mycsreg/CSReg[2][18] ;
wire \mycsreg/CSReg[2][19] ;
wire \mycsreg/CSReg[2][1] ;
wire \mycsreg/CSReg[2][20] ;
wire \mycsreg/CSReg[2][21] ;
wire \mycsreg/CSReg[2][22] ;
wire \mycsreg/CSReg[2][23] ;
wire \mycsreg/CSReg[2][24] ;
wire \mycsreg/CSReg[2][25] ;
wire \mycsreg/CSReg[2][26] ;
wire \mycsreg/CSReg[2][27] ;
wire \mycsreg/CSReg[2][28] ;
wire \mycsreg/CSReg[2][29] ;
wire \mycsreg/CSReg[2][2] ;
wire \mycsreg/CSReg[2][30] ;
wire \mycsreg/CSReg[2][31] ;
wire \mycsreg/CSReg[2][3] ;
wire \mycsreg/CSReg[2][4] ;
wire \mycsreg/CSReg[2][5] ;
wire \mycsreg/CSReg[2][6] ;
wire \mycsreg/CSReg[2][7] ;
wire \mycsreg/CSReg[2][8] ;
wire \mycsreg/CSReg[2][9] ;
wire \mycsreg/CSReg[3][0] ;
wire \mycsreg/CSReg[3][10] ;
wire \mycsreg/CSReg[3][11] ;
wire \mycsreg/CSReg[3][12] ;
wire \mycsreg/CSReg[3][13] ;
wire \mycsreg/CSReg[3][14] ;
wire \mycsreg/CSReg[3][15] ;
wire \mycsreg/CSReg[3][16] ;
wire \mycsreg/CSReg[3][17] ;
wire \mycsreg/CSReg[3][18] ;
wire \mycsreg/CSReg[3][19] ;
wire \mycsreg/CSReg[3][1] ;
wire \mycsreg/CSReg[3][20] ;
wire \mycsreg/CSReg[3][21] ;
wire \mycsreg/CSReg[3][22] ;
wire \mycsreg/CSReg[3][23] ;
wire \mycsreg/CSReg[3][24] ;
wire \mycsreg/CSReg[3][25] ;
wire \mycsreg/CSReg[3][26] ;
wire \mycsreg/CSReg[3][27] ;
wire \mycsreg/CSReg[3][28] ;
wire \mycsreg/CSReg[3][29] ;
wire \mycsreg/CSReg[3][2] ;
wire \mycsreg/CSReg[3][30] ;
wire \mycsreg/CSReg[3][31] ;
wire \mycsreg/CSReg[3][3] ;
wire \mycsreg/CSReg[3][4] ;
wire \mycsreg/CSReg[3][5] ;
wire \mycsreg/CSReg[3][6] ;
wire \mycsreg/CSReg[3][7] ;
wire \mycsreg/CSReg[3][8] ;
wire \mycsreg/CSReg[3][9] ;
wire \myexu/_0000_ ;
wire \myexu/_0001_ ;
wire \myexu/_0002_ ;
wire \myexu/_0003_ ;
wire \myexu/_0004_ ;
wire \myexu/_0005_ ;
wire \myexu/_0006_ ;
wire \myexu/_0007_ ;
wire \myexu/_0008_ ;
wire \myexu/_0009_ ;
wire \myexu/_0010_ ;
wire \myexu/_0011_ ;
wire \myexu/_0012_ ;
wire \myexu/_0013_ ;
wire \myexu/_0014_ ;
wire \myexu/_0015_ ;
wire \myexu/_0016_ ;
wire \myexu/_0017_ ;
wire \myexu/_0018_ ;
wire \myexu/_0019_ ;
wire \myexu/_0020_ ;
wire \myexu/_0021_ ;
wire \myexu/_0022_ ;
wire \myexu/_0023_ ;
wire \myexu/_0024_ ;
wire \myexu/_0025_ ;
wire \myexu/_0026_ ;
wire \myexu/_0027_ ;
wire \myexu/_0028_ ;
wire \myexu/_0029_ ;
wire \myexu/_0030_ ;
wire \myexu/_0031_ ;
wire \myexu/_0032_ ;
wire \myexu/_0033_ ;
wire \myexu/_0034_ ;
wire \myexu/_0035_ ;
wire \myexu/_0036_ ;
wire \myexu/_0037_ ;
wire \myexu/_0038_ ;
wire \myexu/_0039_ ;
wire \myexu/_0040_ ;
wire \myexu/_0041_ ;
wire \myexu/_0042_ ;
wire \myexu/_0043_ ;
wire \myexu/_0044_ ;
wire \myexu/_0045_ ;
wire \myexu/_0046_ ;
wire \myexu/_0047_ ;
wire \myexu/_0048_ ;
wire \myexu/_0049_ ;
wire \myexu/_0050_ ;
wire \myexu/_0051_ ;
wire \myexu/_0052_ ;
wire \myexu/_0053_ ;
wire \myexu/_0054_ ;
wire \myexu/_0055_ ;
wire \myexu/_0056_ ;
wire \myexu/_0057_ ;
wire \myexu/_0058_ ;
wire \myexu/_0059_ ;
wire \myexu/_0060_ ;
wire \myexu/_0061_ ;
wire \myexu/_0062_ ;
wire \myexu/_0063_ ;
wire \myexu/_0064_ ;
wire \myexu/_0065_ ;
wire \myexu/_0066_ ;
wire \myexu/_0067_ ;
wire \myexu/_0068_ ;
wire \myexu/_0069_ ;
wire \myexu/_0070_ ;
wire \myexu/_0071_ ;
wire \myexu/_0072_ ;
wire \myexu/_0073_ ;
wire \myexu/_0074_ ;
wire \myexu/_0075_ ;
wire \myexu/_0076_ ;
wire \myexu/_0077_ ;
wire \myexu/_0078_ ;
wire \myexu/_0079_ ;
wire \myexu/_0080_ ;
wire \myexu/_0081_ ;
wire \myexu/_0082_ ;
wire \myexu/_0083_ ;
wire \myexu/_0084_ ;
wire \myexu/_0085_ ;
wire \myexu/_0086_ ;
wire \myexu/_0087_ ;
wire \myexu/_0088_ ;
wire \myexu/_0089_ ;
wire \myexu/_0090_ ;
wire \myexu/_0091_ ;
wire \myexu/_0092_ ;
wire \myexu/_0093_ ;
wire \myexu/_0094_ ;
wire \myexu/_0095_ ;
wire \myexu/_0096_ ;
wire \myexu/_0097_ ;
wire \myexu/_0098_ ;
wire \myexu/_0099_ ;
wire \myexu/_0100_ ;
wire \myexu/_0101_ ;
wire \myexu/_0102_ ;
wire \myexu/_0103_ ;
wire \myexu/_0104_ ;
wire \myexu/_0105_ ;
wire \myexu/_0106_ ;
wire \myexu/_0107_ ;
wire \myexu/_0108_ ;
wire \myexu/_0109_ ;
wire \myexu/_0110_ ;
wire \myexu/_0111_ ;
wire \myexu/_0112_ ;
wire \myexu/_0113_ ;
wire \myexu/_0114_ ;
wire \myexu/_0115_ ;
wire \myexu/_0116_ ;
wire \myexu/_0117_ ;
wire \myexu/_0118_ ;
wire \myexu/_0119_ ;
wire \myexu/_0120_ ;
wire \myexu/_0121_ ;
wire \myexu/_0122_ ;
wire \myexu/_0123_ ;
wire \myexu/_0124_ ;
wire \myexu/_0125_ ;
wire \myexu/_0126_ ;
wire \myexu/_0127_ ;
wire \myexu/_0128_ ;
wire \myexu/_0129_ ;
wire \myexu/_0130_ ;
wire \myexu/_0131_ ;
wire \myexu/_0132_ ;
wire \myexu/_0133_ ;
wire \myexu/_0134_ ;
wire \myexu/_0135_ ;
wire \myexu/_0136_ ;
wire \myexu/_0137_ ;
wire \myexu/_0138_ ;
wire \myexu/_0139_ ;
wire \myexu/_0140_ ;
wire \myexu/_0141_ ;
wire \myexu/_0142_ ;
wire \myexu/_0143_ ;
wire \myexu/_0144_ ;
wire \myexu/_0145_ ;
wire \myexu/_0146_ ;
wire \myexu/_0147_ ;
wire \myexu/_0148_ ;
wire \myexu/_0149_ ;
wire \myexu/_0150_ ;
wire \myexu/_0151_ ;
wire \myexu/_0152_ ;
wire \myexu/_0153_ ;
wire \myexu/_0154_ ;
wire \myexu/_0155_ ;
wire \myexu/_0156_ ;
wire \myexu/_0157_ ;
wire \myexu/_0158_ ;
wire \myexu/_0159_ ;
wire \myexu/_0160_ ;
wire \myexu/_0161_ ;
wire \myexu/_0162_ ;
wire \myexu/_0163_ ;
wire \myexu/_0164_ ;
wire \myexu/_0165_ ;
wire \myexu/_0166_ ;
wire \myexu/_0167_ ;
wire \myexu/_0168_ ;
wire \myexu/_0169_ ;
wire \myexu/_0170_ ;
wire \myexu/_0171_ ;
wire \myexu/_0172_ ;
wire \myexu/_0173_ ;
wire \myexu/_0174_ ;
wire \myexu/_0175_ ;
wire \myexu/_0176_ ;
wire \myexu/_0177_ ;
wire \myexu/_0178_ ;
wire \myexu/_0179_ ;
wire \myexu/_0180_ ;
wire \myexu/_0181_ ;
wire \myexu/_0182_ ;
wire \myexu/_0183_ ;
wire \myexu/_0184_ ;
wire \myexu/_0185_ ;
wire \myexu/_0186_ ;
wire \myexu/_0187_ ;
wire \myexu/_0188_ ;
wire \myexu/_0189_ ;
wire \myexu/_0190_ ;
wire \myexu/_0191_ ;
wire \myexu/_0192_ ;
wire \myexu/_0193_ ;
wire \myexu/_0194_ ;
wire \myexu/_0195_ ;
wire \myexu/_0196_ ;
wire \myexu/_0197_ ;
wire \myexu/_0198_ ;
wire \myexu/_0199_ ;
wire \myexu/_0200_ ;
wire \myexu/_0201_ ;
wire \myexu/_0202_ ;
wire \myexu/_0203_ ;
wire \myexu/_0204_ ;
wire \myexu/_0205_ ;
wire \myexu/_0206_ ;
wire \myexu/_0207_ ;
wire \myexu/_0208_ ;
wire \myexu/_0209_ ;
wire \myexu/_0210_ ;
wire \myexu/_0211_ ;
wire \myexu/_0212_ ;
wire \myexu/_0213_ ;
wire \myexu/_0214_ ;
wire \myexu/_0215_ ;
wire \myexu/_0216_ ;
wire \myexu/_0217_ ;
wire \myexu/_0218_ ;
wire \myexu/_0219_ ;
wire \myexu/_0220_ ;
wire \myexu/_0221_ ;
wire \myexu/_0222_ ;
wire \myexu/_0223_ ;
wire \myexu/_0224_ ;
wire \myexu/_0225_ ;
wire \myexu/_0226_ ;
wire \myexu/_0227_ ;
wire \myexu/_0228_ ;
wire \myexu/_0229_ ;
wire \myexu/_0230_ ;
wire \myexu/_0231_ ;
wire \myexu/_0232_ ;
wire \myexu/_0233_ ;
wire \myexu/_0234_ ;
wire \myexu/_0235_ ;
wire \myexu/_0236_ ;
wire \myexu/_0237_ ;
wire \myexu/_0238_ ;
wire \myexu/_0239_ ;
wire \myexu/_0240_ ;
wire \myexu/_0241_ ;
wire \myexu/_0242_ ;
wire \myexu/_0243_ ;
wire \myexu/_0244_ ;
wire \myexu/_0245_ ;
wire \myexu/_0246_ ;
wire \myexu/_0247_ ;
wire \myexu/_0248_ ;
wire \myexu/_0249_ ;
wire \myexu/_0250_ ;
wire \myexu/_0251_ ;
wire \myexu/_0252_ ;
wire \myexu/_0253_ ;
wire \myexu/_0254_ ;
wire \myexu/_0255_ ;
wire \myexu/_0256_ ;
wire \myexu/_0257_ ;
wire \myexu/_0258_ ;
wire \myexu/_0259_ ;
wire \myexu/_0260_ ;
wire \myexu/_0261_ ;
wire \myexu/_0262_ ;
wire \myexu/_0263_ ;
wire \myexu/_0264_ ;
wire \myexu/_0265_ ;
wire \myexu/_0266_ ;
wire \myexu/_0267_ ;
wire \myexu/_0268_ ;
wire \myexu/_0269_ ;
wire \myexu/_0270_ ;
wire \myexu/_0271_ ;
wire \myexu/_0272_ ;
wire \myexu/_0273_ ;
wire \myexu/_0274_ ;
wire \myexu/_0275_ ;
wire \myexu/_0276_ ;
wire \myexu/_0277_ ;
wire \myexu/_0278_ ;
wire \myexu/_0279_ ;
wire \myexu/_0280_ ;
wire \myexu/_0281_ ;
wire \myexu/_0282_ ;
wire \myexu/_0283_ ;
wire \myexu/_0284_ ;
wire \myexu/_0285_ ;
wire \myexu/_0286_ ;
wire \myexu/_0287_ ;
wire \myexu/_0288_ ;
wire \myexu/_0289_ ;
wire \myexu/_0290_ ;
wire \myexu/_0291_ ;
wire \myexu/_0292_ ;
wire \myexu/_0293_ ;
wire \myexu/_0294_ ;
wire \myexu/_0295_ ;
wire \myexu/_0296_ ;
wire \myexu/_0297_ ;
wire \myexu/_0298_ ;
wire \myexu/_0299_ ;
wire \myexu/_0300_ ;
wire \myexu/_0301_ ;
wire \myexu/_0302_ ;
wire \myexu/_0303_ ;
wire \myexu/_0304_ ;
wire \myexu/_0305_ ;
wire \myexu/_0306_ ;
wire \myexu/_0307_ ;
wire \myexu/_0308_ ;
wire \myexu/_0309_ ;
wire \myexu/_0310_ ;
wire \myexu/_0311_ ;
wire \myexu/_0312_ ;
wire \myexu/_0313_ ;
wire \myexu/_0314_ ;
wire \myexu/_0315_ ;
wire \myexu/_0316_ ;
wire \myexu/_0317_ ;
wire \myexu/_0318_ ;
wire \myexu/_0319_ ;
wire \myexu/_0320_ ;
wire \myexu/_0321_ ;
wire \myexu/_0322_ ;
wire \myexu/_0323_ ;
wire \myexu/_0324_ ;
wire \myexu/_0325_ ;
wire \myexu/_0326_ ;
wire \myexu/_0327_ ;
wire \myexu/_0328_ ;
wire \myexu/_0329_ ;
wire \myexu/_0330_ ;
wire \myexu/_0331_ ;
wire \myexu/_0332_ ;
wire \myexu/_0333_ ;
wire \myexu/_0334_ ;
wire \myexu/_0335_ ;
wire \myexu/_0336_ ;
wire \myexu/_0337_ ;
wire \myexu/_0338_ ;
wire \myexu/_0339_ ;
wire \myexu/_0340_ ;
wire \myexu/_0341_ ;
wire \myexu/_0342_ ;
wire \myexu/_0343_ ;
wire \myexu/_0344_ ;
wire \myexu/_0345_ ;
wire \myexu/_0346_ ;
wire \myexu/_0347_ ;
wire \myexu/_0348_ ;
wire \myexu/_0349_ ;
wire \myexu/_0350_ ;
wire \myexu/_0351_ ;
wire \myexu/_0352_ ;
wire \myexu/_0353_ ;
wire \myexu/_0354_ ;
wire \myexu/_0355_ ;
wire \myexu/_0356_ ;
wire \myexu/_0357_ ;
wire \myexu/_0358_ ;
wire \myexu/_0359_ ;
wire \myexu/_0360_ ;
wire \myexu/_0361_ ;
wire \myexu/_0362_ ;
wire \myexu/_0363_ ;
wire \myexu/_0364_ ;
wire \myexu/_0365_ ;
wire \myexu/_0366_ ;
wire \myexu/_0367_ ;
wire \myexu/_0368_ ;
wire \myexu/_0369_ ;
wire \myexu/_0370_ ;
wire \myexu/_0371_ ;
wire \myexu/_0372_ ;
wire \myexu/_0373_ ;
wire \myexu/_0374_ ;
wire \myexu/_0375_ ;
wire \myexu/_0376_ ;
wire \myexu/_0377_ ;
wire \myexu/_0378_ ;
wire \myexu/_0379_ ;
wire \myexu/_0380_ ;
wire \myexu/_0381_ ;
wire \myexu/_0382_ ;
wire \myexu/_0383_ ;
wire \myexu/_0384_ ;
wire \myexu/_0385_ ;
wire \myexu/_0386_ ;
wire \myexu/_0387_ ;
wire \myexu/_0388_ ;
wire \myexu/_0389_ ;
wire \myexu/_0390_ ;
wire \myexu/_0391_ ;
wire \myexu/_0392_ ;
wire \myexu/_0393_ ;
wire \myexu/_0394_ ;
wire \myexu/_0395_ ;
wire \myexu/_0396_ ;
wire \myexu/_0397_ ;
wire \myexu/_0398_ ;
wire \myexu/_0399_ ;
wire \myexu/_0400_ ;
wire \myexu/_0401_ ;
wire \myexu/_0402_ ;
wire \myexu/_0403_ ;
wire \myexu/_0404_ ;
wire \myexu/_0405_ ;
wire \myexu/_0406_ ;
wire \myexu/_0407_ ;
wire \myexu/_0408_ ;
wire \myexu/_0409_ ;
wire \myexu/_0410_ ;
wire \myexu/_0411_ ;
wire \myexu/_0412_ ;
wire \myexu/_0413_ ;
wire \myexu/_0414_ ;
wire \myexu/_0415_ ;
wire \myexu/_0416_ ;
wire \myexu/_0417_ ;
wire \myexu/_0418_ ;
wire \myexu/_0419_ ;
wire \myexu/_0420_ ;
wire \myexu/_0421_ ;
wire \myexu/_0422_ ;
wire \myexu/_0423_ ;
wire \myexu/_0424_ ;
wire \myexu/_0425_ ;
wire \myexu/_0426_ ;
wire \myexu/_0427_ ;
wire \myexu/_0428_ ;
wire \myexu/_0429_ ;
wire \myexu/_0430_ ;
wire \myexu/_0431_ ;
wire \myexu/_0432_ ;
wire \myexu/_0433_ ;
wire \myexu/_0434_ ;
wire \myexu/_0435_ ;
wire \myexu/_0436_ ;
wire \myexu/_0437_ ;
wire \myexu/_0438_ ;
wire \myexu/_0439_ ;
wire \myexu/_0440_ ;
wire \myexu/_0441_ ;
wire \myexu/_0442_ ;
wire \myexu/_0443_ ;
wire \myexu/_0444_ ;
wire \myexu/_0445_ ;
wire \myexu/_0446_ ;
wire \myexu/_0447_ ;
wire \myexu/_0448_ ;
wire \myexu/_0449_ ;
wire \myexu/_0450_ ;
wire \myexu/_0451_ ;
wire \myexu/_0452_ ;
wire \myexu/_0453_ ;
wire \myexu/_0454_ ;
wire \myexu/_0455_ ;
wire \myexu/_0456_ ;
wire \myexu/_0457_ ;
wire \myexu/_0458_ ;
wire \myexu/_0459_ ;
wire \myexu/_0460_ ;
wire \myexu/_0461_ ;
wire \myexu/_0462_ ;
wire \myexu/_0463_ ;
wire \myexu/_0464_ ;
wire \myexu/_0465_ ;
wire \myexu/_0466_ ;
wire \myexu/_0467_ ;
wire \myexu/_0468_ ;
wire \myexu/_0469_ ;
wire \myexu/_0470_ ;
wire \myexu/_0471_ ;
wire \myexu/_0472_ ;
wire \myexu/_0473_ ;
wire \myexu/_0474_ ;
wire \myexu/_0475_ ;
wire \myexu/_0476_ ;
wire \myexu/_0477_ ;
wire \myexu/_0478_ ;
wire \myexu/_0479_ ;
wire \myexu/_0480_ ;
wire \myexu/_0481_ ;
wire \myexu/_0482_ ;
wire \myexu/_0483_ ;
wire \myexu/_0484_ ;
wire \myexu/_0485_ ;
wire \myexu/_0486_ ;
wire \myexu/_0487_ ;
wire \myexu/_0488_ ;
wire \myexu/_0489_ ;
wire \myexu/_0490_ ;
wire \myexu/_0491_ ;
wire \myexu/_0492_ ;
wire \myexu/_0493_ ;
wire \myexu/_0494_ ;
wire \myexu/_0495_ ;
wire \myexu/_0496_ ;
wire \myexu/_0497_ ;
wire \myexu/_0498_ ;
wire \myexu/_0499_ ;
wire \myexu/_0500_ ;
wire \myexu/_0501_ ;
wire \myexu/_0502_ ;
wire \myexu/_0503_ ;
wire \myexu/_0504_ ;
wire \myexu/_0505_ ;
wire \myexu/_0506_ ;
wire \myexu/_0507_ ;
wire \myexu/_0508_ ;
wire \myexu/_0509_ ;
wire \myexu/_0510_ ;
wire \myexu/_0511_ ;
wire \myexu/_0512_ ;
wire \myexu/_0513_ ;
wire \myexu/_0514_ ;
wire \myexu/_0515_ ;
wire \myexu/_0516_ ;
wire \myexu/_0517_ ;
wire \myexu/_0518_ ;
wire \myexu/_0519_ ;
wire \myexu/_0520_ ;
wire \myexu/_0521_ ;
wire \myexu/_0522_ ;
wire \myexu/_0523_ ;
wire \myexu/_0524_ ;
wire \myexu/_0525_ ;
wire \myexu/_0526_ ;
wire \myexu/_0527_ ;
wire \myexu/_0528_ ;
wire \myexu/_0529_ ;
wire \myexu/_0530_ ;
wire \myexu/_0531_ ;
wire \myexu/_0532_ ;
wire \myexu/_0533_ ;
wire \myexu/_0534_ ;
wire \myexu/_0535_ ;
wire \myexu/_0536_ ;
wire \myexu/_0537_ ;
wire \myexu/_0538_ ;
wire \myexu/_0539_ ;
wire \myexu/_0540_ ;
wire \myexu/_0541_ ;
wire \myexu/_0542_ ;
wire \myexu/_0543_ ;
wire \myexu/_0544_ ;
wire \myexu/_0545_ ;
wire \myexu/_0546_ ;
wire \myexu/_0547_ ;
wire \myexu/_0548_ ;
wire \myexu/_0549_ ;
wire \myexu/_0550_ ;
wire \myexu/_0551_ ;
wire \myexu/_0552_ ;
wire \myexu/_0553_ ;
wire \myexu/_0554_ ;
wire \myexu/_0555_ ;
wire \myexu/_0556_ ;
wire \myexu/_0557_ ;
wire \myexu/_0558_ ;
wire \myexu/_0559_ ;
wire \myexu/_0560_ ;
wire \myexu/_0561_ ;
wire \myexu/_0562_ ;
wire \myexu/_0563_ ;
wire \myexu/_0564_ ;
wire \myexu/_0565_ ;
wire \myexu/_0566_ ;
wire \myexu/_0567_ ;
wire \myexu/_0568_ ;
wire \myexu/_0569_ ;
wire \myexu/_0570_ ;
wire \myexu/_0571_ ;
wire \myexu/_0572_ ;
wire \myexu/_0573_ ;
wire \myexu/_0574_ ;
wire \myexu/_0575_ ;
wire \myexu/_0576_ ;
wire \myexu/_0577_ ;
wire \myexu/_0578_ ;
wire \myexu/_0579_ ;
wire \myexu/_0580_ ;
wire \myexu/_0581_ ;
wire \myexu/_0582_ ;
wire \myexu/_0583_ ;
wire \myexu/_0584_ ;
wire \myexu/_0585_ ;
wire \myexu/_0586_ ;
wire \myexu/_0587_ ;
wire \myexu/_0588_ ;
wire \myexu/_0589_ ;
wire \myexu/_0590_ ;
wire \myexu/_0591_ ;
wire \myexu/_0592_ ;
wire \myexu/_0593_ ;
wire \myexu/_0594_ ;
wire \myexu/_0595_ ;
wire \myexu/_0596_ ;
wire \myexu/_0597_ ;
wire \myexu/_0598_ ;
wire \myexu/_0599_ ;
wire \myexu/_0600_ ;
wire \myexu/_0601_ ;
wire \myexu/_0602_ ;
wire \myexu/_0603_ ;
wire \myexu/_0604_ ;
wire \myexu/_0605_ ;
wire \myexu/_0606_ ;
wire \myexu/_0607_ ;
wire \myexu/_0608_ ;
wire \myexu/_0609_ ;
wire \myexu/_0610_ ;
wire \myexu/_0611_ ;
wire \myexu/_0612_ ;
wire \myexu/_0613_ ;
wire \myexu/_0614_ ;
wire \myexu/_0615_ ;
wire \myexu/_0616_ ;
wire \myexu/_0617_ ;
wire \myexu/_0618_ ;
wire \myexu/_0619_ ;
wire \myexu/_0620_ ;
wire \myexu/_0621_ ;
wire \myexu/_0622_ ;
wire \myexu/_0623_ ;
wire \myexu/_0624_ ;
wire \myexu/_0625_ ;
wire \myexu/_0626_ ;
wire \myexu/_0627_ ;
wire \myexu/_0628_ ;
wire \myexu/_0629_ ;
wire \myexu/_0630_ ;
wire \myexu/_0631_ ;
wire \myexu/_0632_ ;
wire \myexu/_0633_ ;
wire \myexu/_0634_ ;
wire \myexu/_0635_ ;
wire \myexu/_0636_ ;
wire \myexu/_0637_ ;
wire \myexu/_0638_ ;
wire \myexu/_0639_ ;
wire \myexu/_0640_ ;
wire \myexu/_0641_ ;
wire \myexu/_0642_ ;
wire \myexu/_0643_ ;
wire \myexu/_0644_ ;
wire \myexu/_0645_ ;
wire \myexu/_0646_ ;
wire \myexu/_0647_ ;
wire \myexu/_0648_ ;
wire \myexu/_0649_ ;
wire \myexu/_0650_ ;
wire \myexu/_0651_ ;
wire \myexu/_0652_ ;
wire \myexu/_0653_ ;
wire \myexu/_0654_ ;
wire \myexu/_0655_ ;
wire \myexu/_0656_ ;
wire \myexu/_0657_ ;
wire \myexu/_0658_ ;
wire \myexu/_0659_ ;
wire \myexu/_0660_ ;
wire \myexu/_0661_ ;
wire \myexu/_0662_ ;
wire \myexu/_0663_ ;
wire \myexu/_0664_ ;
wire \myexu/_0665_ ;
wire \myexu/_0666_ ;
wire \myexu/_0667_ ;
wire \myexu/_0668_ ;
wire \myexu/_0669_ ;
wire \myexu/_0670_ ;
wire \myexu/_0671_ ;
wire \myexu/_0672_ ;
wire \myexu/_0673_ ;
wire \myexu/_0674_ ;
wire \myexu/_0675_ ;
wire \myexu/_0676_ ;
wire \myexu/_0677_ ;
wire \myexu/_0678_ ;
wire \myexu/_0679_ ;
wire \myexu/_0680_ ;
wire \myexu/_0681_ ;
wire \myexu/_0682_ ;
wire \myexu/_0683_ ;
wire \myexu/_0684_ ;
wire \myexu/_0685_ ;
wire \myexu/_0686_ ;
wire \myexu/_0687_ ;
wire \myexu/_0688_ ;
wire \myexu/_0689_ ;
wire \myexu/_0690_ ;
wire \myexu/_0691_ ;
wire \myexu/_0692_ ;
wire \myexu/_0693_ ;
wire \myexu/_0694_ ;
wire \myexu/_0695_ ;
wire \myexu/_0696_ ;
wire \myexu/_0697_ ;
wire \myexu/_0698_ ;
wire \myexu/_0699_ ;
wire \myexu/_0700_ ;
wire \myexu/_0701_ ;
wire \myexu/_0702_ ;
wire \myexu/_0703_ ;
wire \myexu/_0704_ ;
wire \myexu/_0705_ ;
wire \myexu/_0706_ ;
wire \myexu/_0707_ ;
wire \myexu/_0708_ ;
wire \myexu/_0709_ ;
wire \myexu/_0710_ ;
wire \myexu/_0711_ ;
wire \myexu/_0712_ ;
wire \myexu/_0713_ ;
wire \myexu/_0714_ ;
wire \myexu/_0715_ ;
wire \myexu/_0716_ ;
wire \myexu/_0717_ ;
wire \myexu/_0718_ ;
wire \myexu/_0719_ ;
wire \myexu/_0720_ ;
wire \myexu/_0721_ ;
wire \myexu/_0722_ ;
wire \myexu/_0723_ ;
wire \myexu/_0724_ ;
wire \myexu/_0725_ ;
wire \myexu/_0726_ ;
wire \myexu/_0727_ ;
wire \myexu/_0728_ ;
wire \myexu/_0729_ ;
wire \myexu/_0730_ ;
wire \myexu/_0731_ ;
wire \myexu/_0732_ ;
wire \myexu/_0733_ ;
wire \myexu/_0734_ ;
wire \myexu/_0735_ ;
wire \myexu/_0736_ ;
wire \myexu/_0737_ ;
wire \myexu/_0738_ ;
wire \myexu/_0739_ ;
wire \myexu/_0740_ ;
wire \myexu/_0741_ ;
wire \myexu/_0742_ ;
wire \myexu/_0743_ ;
wire \myexu/_0744_ ;
wire \myexu/_0745_ ;
wire \myexu/_0746_ ;
wire \myexu/_0747_ ;
wire \myexu/_0748_ ;
wire \myexu/_0749_ ;
wire \myexu/_0750_ ;
wire \myexu/_0751_ ;
wire \myexu/_0752_ ;
wire \myexu/_0753_ ;
wire \myexu/_0754_ ;
wire \myexu/_0755_ ;
wire \myexu/_0756_ ;
wire \myexu/_0757_ ;
wire \myexu/_0758_ ;
wire \myexu/_0759_ ;
wire \myexu/_0760_ ;
wire \myexu/_0761_ ;
wire \myexu/_0762_ ;
wire \myexu/_0763_ ;
wire \myexu/_0764_ ;
wire \myexu/_0765_ ;
wire \myexu/_0766_ ;
wire \myexu/_0767_ ;
wire \myexu/_0768_ ;
wire \myexu/_0769_ ;
wire \myexu/_0770_ ;
wire \myexu/_0771_ ;
wire \myexu/_0772_ ;
wire \myexu/_0773_ ;
wire \myexu/_0774_ ;
wire \myexu/_0775_ ;
wire \myexu/_0776_ ;
wire \myexu/_0777_ ;
wire \myexu/_0778_ ;
wire \myexu/_0779_ ;
wire \myexu/_0780_ ;
wire \myexu/_0781_ ;
wire \myexu/_0782_ ;
wire \myexu/_0783_ ;
wire \myexu/_0784_ ;
wire \myexu/_0785_ ;
wire \myexu/_0786_ ;
wire \myexu/_0787_ ;
wire \myexu/_0788_ ;
wire \myexu/_0789_ ;
wire \myexu/_0790_ ;
wire \myexu/_0791_ ;
wire \myexu/_0792_ ;
wire \myexu/_0793_ ;
wire \myexu/_0794_ ;
wire \myexu/_0795_ ;
wire \myexu/_0796_ ;
wire \myexu/_0797_ ;
wire \myexu/_0798_ ;
wire \myexu/_0799_ ;
wire \myexu/_0800_ ;
wire \myexu/_0801_ ;
wire \myexu/_0802_ ;
wire \myexu/_0803_ ;
wire \myexu/_0804_ ;
wire \myexu/_0805_ ;
wire \myexu/_0806_ ;
wire \myexu/_0807_ ;
wire \myexu/_0808_ ;
wire \myexu/_0809_ ;
wire \myexu/_0810_ ;
wire \myexu/_0811_ ;
wire \myexu/_0812_ ;
wire \myexu/_0813_ ;
wire \myexu/_0814_ ;
wire \myexu/_0815_ ;
wire \myexu/_0816_ ;
wire \myexu/_0817_ ;
wire \myexu/_0818_ ;
wire \myexu/_0819_ ;
wire \myexu/_0820_ ;
wire \myexu/_0821_ ;
wire \myexu/_0822_ ;
wire \myexu/_0823_ ;
wire \myexu/_0824_ ;
wire \myexu/_0825_ ;
wire \myexu/_0826_ ;
wire \myexu/_0827_ ;
wire \myexu/_0828_ ;
wire \myexu/_0829_ ;
wire \myexu/_0830_ ;
wire \myexu/_0831_ ;
wire \myexu/_0832_ ;
wire \myexu/_0833_ ;
wire \myexu/_0834_ ;
wire \myexu/_0835_ ;
wire \myexu/_0836_ ;
wire \myexu/_0837_ ;
wire \myexu/_0838_ ;
wire \myexu/_0839_ ;
wire \myexu/_0840_ ;
wire \myexu/_0841_ ;
wire \myexu/_0842_ ;
wire \myexu/_0843_ ;
wire \myexu/_0844_ ;
wire \myexu/_0845_ ;
wire \myexu/_0846_ ;
wire \myexu/_0847_ ;
wire \myexu/_0848_ ;
wire \myexu/_0849_ ;
wire \myexu/_0850_ ;
wire \myexu/_0851_ ;
wire \myexu/_0852_ ;
wire \myexu/_0853_ ;
wire \myexu/_0854_ ;
wire \myexu/_0855_ ;
wire \myexu/_0856_ ;
wire \myexu/_0857_ ;
wire \myexu/_0858_ ;
wire \myexu/_0859_ ;
wire \myexu/_0860_ ;
wire \myexu/_0861_ ;
wire \myexu/_0862_ ;
wire \myexu/_0863_ ;
wire \myexu/_0864_ ;
wire \myexu/_0865_ ;
wire \myexu/_0866_ ;
wire \myexu/_0867_ ;
wire \myexu/_0868_ ;
wire \myexu/_0869_ ;
wire \myexu/_0870_ ;
wire \myexu/_0871_ ;
wire \myexu/_0872_ ;
wire \myexu/_0873_ ;
wire \myexu/_0874_ ;
wire \myexu/_0875_ ;
wire \myexu/_0876_ ;
wire \myexu/_0877_ ;
wire \myexu/_0878_ ;
wire \myexu/_0879_ ;
wire \myexu/_0880_ ;
wire \myexu/_0881_ ;
wire \myexu/_0882_ ;
wire \myexu/_0883_ ;
wire \myexu/_0884_ ;
wire \myexu/_0885_ ;
wire \myexu/_0886_ ;
wire \myexu/_0887_ ;
wire \myexu/_0888_ ;
wire \myexu/_0889_ ;
wire \myexu/_0890_ ;
wire \myexu/_0891_ ;
wire \myexu/_0892_ ;
wire \myexu/_0893_ ;
wire \myexu/_0894_ ;
wire \myexu/_0895_ ;
wire \myexu/_0896_ ;
wire \myexu/_0897_ ;
wire \myexu/_0898_ ;
wire \myexu/_0899_ ;
wire \myexu/_0900_ ;
wire \myexu/_0901_ ;
wire \myexu/_0902_ ;
wire \myexu/_0903_ ;
wire \myexu/_0904_ ;
wire \myexu/_0905_ ;
wire \myexu/_0906_ ;
wire \myexu/_0907_ ;
wire \myexu/_0908_ ;
wire \myexu/_0909_ ;
wire \myexu/_0910_ ;
wire \myexu/_0911_ ;
wire \myexu/_0912_ ;
wire \myexu/_0913_ ;
wire \myexu/_0914_ ;
wire \myexu/_0915_ ;
wire \myexu/_0916_ ;
wire \myexu/_0917_ ;
wire \myexu/_0918_ ;
wire \myexu/_0919_ ;
wire \myexu/_0920_ ;
wire \myexu/_0921_ ;
wire \myexu/_0922_ ;
wire \myexu/_0923_ ;
wire \myexu/_0924_ ;
wire \myexu/_0925_ ;
wire \myexu/_0926_ ;
wire \myexu/_0927_ ;
wire \myexu/_0928_ ;
wire \myexu/_0929_ ;
wire \myexu/_0930_ ;
wire \myexu/_0931_ ;
wire \myexu/_0932_ ;
wire \myexu/_0933_ ;
wire \myexu/_0934_ ;
wire \myexu/_0935_ ;
wire \myexu/_0936_ ;
wire \myexu/_0937_ ;
wire \myexu/_0938_ ;
wire \myexu/_0939_ ;
wire \myexu/_0940_ ;
wire \myexu/_0941_ ;
wire \myexu/_0942_ ;
wire \myexu/_0943_ ;
wire \myexu/_0944_ ;
wire \myexu/_0945_ ;
wire \myexu/_0946_ ;
wire \myexu/_0947_ ;
wire \myexu/_0948_ ;
wire \myexu/_0949_ ;
wire \myexu/_0950_ ;
wire \myexu/_0951_ ;
wire \myexu/_0952_ ;
wire \myexu/_0953_ ;
wire \myexu/_0954_ ;
wire \myexu/_0955_ ;
wire \myexu/_0956_ ;
wire \myexu/_0957_ ;
wire \myexu/_0958_ ;
wire \myexu/_0959_ ;
wire \myexu/_0960_ ;
wire \myexu/_0961_ ;
wire \myexu/_0962_ ;
wire \myexu/_0963_ ;
wire \myexu/_0964_ ;
wire \myexu/_0965_ ;
wire \myexu/_0966_ ;
wire \myexu/_0967_ ;
wire \myexu/_0968_ ;
wire \myexu/_0969_ ;
wire \myexu/_0970_ ;
wire \myexu/_0971_ ;
wire \myexu/_0972_ ;
wire \myexu/_0973_ ;
wire \myexu/_0974_ ;
wire \myexu/_0975_ ;
wire \myexu/_0976_ ;
wire \myexu/_0977_ ;
wire \myexu/_0978_ ;
wire \myexu/_0979_ ;
wire \myexu/_0980_ ;
wire \myexu/_0981_ ;
wire \myexu/_0982_ ;
wire \myexu/_0983_ ;
wire \myexu/_0984_ ;
wire \myexu/_0985_ ;
wire \myexu/_0986_ ;
wire \myexu/_0987_ ;
wire \myexu/_0988_ ;
wire \myexu/_0989_ ;
wire \myexu/_0990_ ;
wire \myexu/_0991_ ;
wire \myexu/_0992_ ;
wire \myexu/_0993_ ;
wire \myexu/_0994_ ;
wire \myexu/_0995_ ;
wire \myexu/_0996_ ;
wire \myexu/_0997_ ;
wire \myexu/_0998_ ;
wire \myexu/_0999_ ;
wire \myexu/_1000_ ;
wire \myexu/_1001_ ;
wire \myexu/_1002_ ;
wire \myexu/_1003_ ;
wire \myexu/_1004_ ;
wire \myexu/_1005_ ;
wire \myexu/_1006_ ;
wire \myexu/_1007_ ;
wire \myexu/_1008_ ;
wire \myexu/_1009_ ;
wire \myexu/_1010_ ;
wire \myexu/_1011_ ;
wire \myexu/_1012_ ;
wire \myexu/_1013_ ;
wire \myexu/_1014_ ;
wire \myexu/_1015_ ;
wire \myexu/_1016_ ;
wire \myexu/_1017_ ;
wire \myexu/_1018_ ;
wire \myexu/_1019_ ;
wire \myexu/_1020_ ;
wire \myexu/_1021_ ;
wire \myexu/_1022_ ;
wire \myexu/_1023_ ;
wire \myexu/_1024_ ;
wire \myexu/_1025_ ;
wire \myexu/_1026_ ;
wire \myexu/_1027_ ;
wire \myexu/_1028_ ;
wire \myexu/_1029_ ;
wire \myexu/_1030_ ;
wire \myexu/_1031_ ;
wire \myexu/_1032_ ;
wire \myexu/_1033_ ;
wire \myexu/_1034_ ;
wire \myexu/_1035_ ;
wire \myexu/_1036_ ;
wire \myexu/_1037_ ;
wire \myexu/_1038_ ;
wire \myexu/_1039_ ;
wire \myexu/_1040_ ;
wire \myexu/_1041_ ;
wire \myexu/_1042_ ;
wire \myexu/_1043_ ;
wire \myexu/_1044_ ;
wire \myexu/_1045_ ;
wire \myexu/_1046_ ;
wire \myexu/_1047_ ;
wire \myexu/_1048_ ;
wire \myexu/_1049_ ;
wire \myexu/_1050_ ;
wire \myexu/_1051_ ;
wire \myexu/_1052_ ;
wire \myexu/_1053_ ;
wire \myexu/_1054_ ;
wire \myexu/_1055_ ;
wire \myexu/_1056_ ;
wire \myexu/_1057_ ;
wire \myexu/_1058_ ;
wire \myexu/_1059_ ;
wire \myexu/_1060_ ;
wire \myexu/_1061_ ;
wire \myexu/_1062_ ;
wire \myexu/_1063_ ;
wire \myexu/_1064_ ;
wire \myexu/_1065_ ;
wire \myexu/_1066_ ;
wire \myexu/_1067_ ;
wire \myexu/_1068_ ;
wire \myexu/_1069_ ;
wire \myexu/_1070_ ;
wire \myexu/_1071_ ;
wire \myexu/_1072_ ;
wire \myexu/_1073_ ;
wire \myexu/_1074_ ;
wire \myexu/_1075_ ;
wire \myexu/_1076_ ;
wire \myexu/_1077_ ;
wire \myexu/_1078_ ;
wire \myexu/_1079_ ;
wire \myexu/_1080_ ;
wire \myexu/_1081_ ;
wire \myexu/_1082_ ;
wire \myexu/_1083_ ;
wire \myexu/_1084_ ;
wire \myexu/_1085_ ;
wire \myexu/_1086_ ;
wire \myexu/_1087_ ;
wire \myexu/_1088_ ;
wire \myexu/_1089_ ;
wire \myexu/_1090_ ;
wire \myexu/_1091_ ;
wire \myexu/_1092_ ;
wire \myexu/_1093_ ;
wire \myexu/_1094_ ;
wire \myexu/_1095_ ;
wire \myexu/_1096_ ;
wire \myexu/_1097_ ;
wire \myexu/_1098_ ;
wire \myexu/_1099_ ;
wire \myexu/_1100_ ;
wire \myexu/_1101_ ;
wire \myexu/_1102_ ;
wire \myexu/_1103_ ;
wire \myexu/_1104_ ;
wire \myexu/_1105_ ;
wire \myexu/_1106_ ;
wire \myexu/_1107_ ;
wire \myexu/_1108_ ;
wire \myexu/_1109_ ;
wire \myexu/_1110_ ;
wire \myexu/_1111_ ;
wire \myexu/_1112_ ;
wire \myexu/_1113_ ;
wire \myexu/_1114_ ;
wire \myexu/_1115_ ;
wire \myexu/_1116_ ;
wire \myexu/_1117_ ;
wire \myexu/_1118_ ;
wire \myexu/_1119_ ;
wire \myexu/_1120_ ;
wire \myexu/_1121_ ;
wire \myexu/_1122_ ;
wire \myexu/_1123_ ;
wire \myexu/_1124_ ;
wire \myexu/_1125_ ;
wire \myexu/_1126_ ;
wire \myexu/_1127_ ;
wire \myexu/_1128_ ;
wire \myexu/_1129_ ;
wire \myexu/_1130_ ;
wire \myexu/_1131_ ;
wire \myexu/_1132_ ;
wire \myexu/_1133_ ;
wire \myexu/_1134_ ;
wire \myexu/_1135_ ;
wire \myexu/_1136_ ;
wire \myexu/_1137_ ;
wire \myexu/_1138_ ;
wire \myexu/_1139_ ;
wire \myexu/_1140_ ;
wire \myexu/_1141_ ;
wire \myexu/_1142_ ;
wire \myexu/_1143_ ;
wire \myexu/_1144_ ;
wire \myexu/_1145_ ;
wire \myexu/_1146_ ;
wire \myexu/_1147_ ;
wire \myexu/_1148_ ;
wire \myexu/_1149_ ;
wire \myexu/_1150_ ;
wire \myexu/_1151_ ;
wire \myexu/_1152_ ;
wire \myexu/_1153_ ;
wire \myexu/_1154_ ;
wire \myexu/_1155_ ;
wire \myexu/_1156_ ;
wire \myexu/_1157_ ;
wire \myexu/_1158_ ;
wire \myexu/_1159_ ;
wire \myexu/_1160_ ;
wire \myexu/_1161_ ;
wire \myexu/_1162_ ;
wire \myexu/_1163_ ;
wire \myexu/_1164_ ;
wire \myexu/_1165_ ;
wire \myexu/_1166_ ;
wire \myexu/_1167_ ;
wire \myexu/_1168_ ;
wire \myexu/_1169_ ;
wire \myexu/_1170_ ;
wire \myexu/_1171_ ;
wire \myexu/_1172_ ;
wire \myexu/_1173_ ;
wire \myexu/_1174_ ;
wire \myexu/_1175_ ;
wire \myexu/_1176_ ;
wire \myexu/_1177_ ;
wire \myexu/_1178_ ;
wire \myexu/_1179_ ;
wire \myexu/_1180_ ;
wire \myexu/_1181_ ;
wire \myexu/_1182_ ;
wire \myexu/_1183_ ;
wire \myexu/_1184_ ;
wire \myexu/_1185_ ;
wire \myexu/_1186_ ;
wire \myexu/_1187_ ;
wire \myexu/_1188_ ;
wire \myexu/_1189_ ;
wire \myexu/_1190_ ;
wire \myexu/_1191_ ;
wire \myexu/_1192_ ;
wire \myexu/_1193_ ;
wire \myexu/_1194_ ;
wire \myexu/_1195_ ;
wire \myexu/_1196_ ;
wire \myexu/_1197_ ;
wire \myexu/_1198_ ;
wire \myexu/_1199_ ;
wire \myexu/_1200_ ;
wire \myexu/_1201_ ;
wire \myexu/_1202_ ;
wire \myexu/_1203_ ;
wire \myexu/_1204_ ;
wire \myexu/_1205_ ;
wire \myexu/_1206_ ;
wire \myexu/_1207_ ;
wire \myexu/_1208_ ;
wire \myexu/_1209_ ;
wire \myexu/_1210_ ;
wire \myexu/_1211_ ;
wire \myexu/_1212_ ;
wire \myexu/_1213_ ;
wire \myexu/_1214_ ;
wire \myexu/_1215_ ;
wire \myexu/_1216_ ;
wire \myexu/_1217_ ;
wire \myexu/_1218_ ;
wire \myexu/_1219_ ;
wire \myexu/_1220_ ;
wire \myexu/_1221_ ;
wire \myexu/_1222_ ;
wire \myexu/_1223_ ;
wire \myexu/_1224_ ;
wire \myexu/_1225_ ;
wire \myexu/_1226_ ;
wire \myexu/_1227_ ;
wire \myexu/_1228_ ;
wire \myexu/_1229_ ;
wire \myexu/_1230_ ;
wire \myexu/_1231_ ;
wire \myexu/_1232_ ;
wire \myexu/_1233_ ;
wire \myexu/_1234_ ;
wire \myexu/_1235_ ;
wire \myexu/_1236_ ;
wire \myexu/_1237_ ;
wire \myexu/_1238_ ;
wire \myexu/_1239_ ;
wire \myexu/_1240_ ;
wire \myexu/_1241_ ;
wire \myexu/_1242_ ;
wire \myexu/_1243_ ;
wire \myexu/_1244_ ;
wire \myexu/_1245_ ;
wire \myexu/_1246_ ;
wire \myexu/_1247_ ;
wire \myexu/_1248_ ;
wire \myexu/_1249_ ;
wire \myexu/_1250_ ;
wire \myexu/_1251_ ;
wire \myexu/_1252_ ;
wire \myexu/_1253_ ;
wire \myexu/_1254_ ;
wire \myexu/_1255_ ;
wire \myexu/_1256_ ;
wire \myexu/_1257_ ;
wire \myexu/_1258_ ;
wire \myexu/_1259_ ;
wire \myexu/_1260_ ;
wire \myexu/_1261_ ;
wire \myexu/_1262_ ;
wire \myexu/_1263_ ;
wire \myexu/_1264_ ;
wire \myexu/_1265_ ;
wire \myexu/_1266_ ;
wire \myexu/_1267_ ;
wire \myexu/_1268_ ;
wire \myexu/_1269_ ;
wire \myexu/_1270_ ;
wire \myexu/_1271_ ;
wire \myexu/_1272_ ;
wire \myexu/_1273_ ;
wire \myexu/_1274_ ;
wire \myexu/_1275_ ;
wire \myexu/_1276_ ;
wire \myexu/_1277_ ;
wire \myexu/_1278_ ;
wire \myexu/_1279_ ;
wire \myexu/_1280_ ;
wire \myexu/_1281_ ;
wire \myexu/_1282_ ;
wire \myexu/_1283_ ;
wire \myexu/_1284_ ;
wire \myexu/_1285_ ;
wire \myexu/_1286_ ;
wire \myexu/_1287_ ;
wire \myexu/_1288_ ;
wire \myexu/_1289_ ;
wire \myexu/_1290_ ;
wire \myexu/_1291_ ;
wire \myexu/_1292_ ;
wire \myexu/_1293_ ;
wire \myexu/_1294_ ;
wire \myexu/_1295_ ;
wire \myexu/_1296_ ;
wire \myexu/_1297_ ;
wire \myexu/_1298_ ;
wire \myexu/_1299_ ;
wire \myexu/_1300_ ;
wire \myexu/_1301_ ;
wire \myexu/_1302_ ;
wire \myexu/_1303_ ;
wire \myexu/_1304_ ;
wire \myexu/_1305_ ;
wire \myexu/_1306_ ;
wire \myexu/_1307_ ;
wire \myexu/_1308_ ;
wire \myexu/_1309_ ;
wire \myexu/_1310_ ;
wire \myexu/_1311_ ;
wire \myexu/_1312_ ;
wire \myexu/_1313_ ;
wire \myexu/_1314_ ;
wire \myexu/_1315_ ;
wire \myexu/_1316_ ;
wire \myexu/_1317_ ;
wire \myexu/_1318_ ;
wire \myexu/_1319_ ;
wire \myexu/_1320_ ;
wire \myexu/_1321_ ;
wire \myexu/_1322_ ;
wire \myexu/_1323_ ;
wire \myexu/_1324_ ;
wire \myexu/_1325_ ;
wire \myexu/_1326_ ;
wire \myexu/_1327_ ;
wire \myexu/_1328_ ;
wire \myexu/_1329_ ;
wire \myexu/_1330_ ;
wire \myexu/_1331_ ;
wire \myexu/_1332_ ;
wire \myexu/_1333_ ;
wire \myexu/_1334_ ;
wire \myexu/_1335_ ;
wire \myexu/_1336_ ;
wire \myexu/_1337_ ;
wire \myexu/_1338_ ;
wire \myexu/_1339_ ;
wire \myexu/_1340_ ;
wire \myexu/_1341_ ;
wire \myexu/_1342_ ;
wire \myexu/_1343_ ;
wire \myexu/_1344_ ;
wire \myexu/_1345_ ;
wire \myexu/_1346_ ;
wire \myexu/_1347_ ;
wire \myexu/_1348_ ;
wire \myexu/_1349_ ;
wire \myexu/_1350_ ;
wire \myexu/_1351_ ;
wire \myexu/_1352_ ;
wire \myexu/_1353_ ;
wire \myexu/_1354_ ;
wire \myexu/_1355_ ;
wire \myexu/_1356_ ;
wire \myexu/_1357_ ;
wire \myexu/_1358_ ;
wire \myexu/_1359_ ;
wire \myexu/_1360_ ;
wire \myexu/_1361_ ;
wire \myexu/_1362_ ;
wire \myexu/_1363_ ;
wire \myexu/_1364_ ;
wire \myexu/_1365_ ;
wire \myexu/_1366_ ;
wire \myexu/_1367_ ;
wire \myexu/_1368_ ;
wire \myexu/_1369_ ;
wire \myexu/_1370_ ;
wire \myexu/_1371_ ;
wire \myexu/_1372_ ;
wire \myexu/_1373_ ;
wire \myexu/_1374_ ;
wire \myexu/_1375_ ;
wire \myexu/_1376_ ;
wire \myexu/_1377_ ;
wire \myexu/_1378_ ;
wire \myexu/_1379_ ;
wire \myexu/_1380_ ;
wire \myexu/_1381_ ;
wire \myexu/_1382_ ;
wire \myexu/_1383_ ;
wire \myexu/_1384_ ;
wire \myexu/_1385_ ;
wire \myexu/_1386_ ;
wire \myexu/_1387_ ;
wire \myexu/_1388_ ;
wire \myexu/_1389_ ;
wire \myexu/_1390_ ;
wire \myexu/_1391_ ;
wire \myexu/_1392_ ;
wire \myexu/_1393_ ;
wire \myexu/_1394_ ;
wire \myexu/_1395_ ;
wire \myexu/_1396_ ;
wire \myexu/_1397_ ;
wire \myexu/_1398_ ;
wire \myexu/_1399_ ;
wire \myexu/_1400_ ;
wire \myexu/_1401_ ;
wire \myexu/_1402_ ;
wire \myexu/_1403_ ;
wire \myexu/_1404_ ;
wire \myexu/_1405_ ;
wire \myexu/_1406_ ;
wire \myexu/_1407_ ;
wire \myexu/_1408_ ;
wire \myexu/_1409_ ;
wire \myexu/_1410_ ;
wire \myexu/_1411_ ;
wire \myexu/_1412_ ;
wire \myexu/_1413_ ;
wire \myexu/_1414_ ;
wire \myexu/_1415_ ;
wire \myexu/_1416_ ;
wire \myexu/_1417_ ;
wire \myexu/_1418_ ;
wire \myexu/_1419_ ;
wire \myexu/_1420_ ;
wire \myexu/_1421_ ;
wire \myexu/_1422_ ;
wire \myexu/_1423_ ;
wire \myexu/_1424_ ;
wire \myexu/_1425_ ;
wire \myexu/_1426_ ;
wire \myexu/_1427_ ;
wire \myexu/_1428_ ;
wire \myexu/_1429_ ;
wire \myexu/_1430_ ;
wire \myexu/_1431_ ;
wire \myexu/_1432_ ;
wire \myexu/_1433_ ;
wire \myexu/_1434_ ;
wire \myexu/_1435_ ;
wire \myexu/_1436_ ;
wire \myexu/_1437_ ;
wire \myexu/_1438_ ;
wire \myexu/_1439_ ;
wire \myexu/_1440_ ;
wire \myexu/_1441_ ;
wire \myexu/_1442_ ;
wire \myexu/_1443_ ;
wire \myexu/_1444_ ;
wire \myexu/_1445_ ;
wire \myexu/_1446_ ;
wire \myexu/_1447_ ;
wire \myexu/_1448_ ;
wire \myexu/_1449_ ;
wire \myexu/_1450_ ;
wire \myexu/_1451_ ;
wire \myexu/_1452_ ;
wire \myexu/_1453_ ;
wire \myexu/_1454_ ;
wire \myexu/_1455_ ;
wire \myexu/_1456_ ;
wire \myexu/_1457_ ;
wire \myexu/_1458_ ;
wire \myexu/_1459_ ;
wire \myexu/_1460_ ;
wire \myexu/_1461_ ;
wire \myexu/_1462_ ;
wire \myexu/_1463_ ;
wire \myexu/_1464_ ;
wire \myexu/_1465_ ;
wire \myexu/_1466_ ;
wire \myexu/_1467_ ;
wire \myexu/_1468_ ;
wire \myexu/_1469_ ;
wire \myexu/_1470_ ;
wire \myexu/_1471_ ;
wire \myexu/_1472_ ;
wire \myexu/_1473_ ;
wire \myexu/_1474_ ;
wire \myexu/_1475_ ;
wire \myexu/_1476_ ;
wire \myexu/_1477_ ;
wire \myexu/_1478_ ;
wire \myexu/_1479_ ;
wire \myexu/_1480_ ;
wire \myexu/_1481_ ;
wire \myexu/_1482_ ;
wire \myexu/_1483_ ;
wire \myexu/_1484_ ;
wire \myexu/_1485_ ;
wire \myexu/_1486_ ;
wire \myexu/_1487_ ;
wire \myexu/_1488_ ;
wire \myexu/_1489_ ;
wire \myexu/_1490_ ;
wire \myexu/_1491_ ;
wire \myexu/_1492_ ;
wire \myexu/_1493_ ;
wire \myexu/_1494_ ;
wire \myexu/_1495_ ;
wire \myexu/_1496_ ;
wire \myexu/_1497_ ;
wire \myexu/_1498_ ;
wire \myexu/_1499_ ;
wire \myexu/_1500_ ;
wire \myexu/_1501_ ;
wire \myexu/_1502_ ;
wire \myexu/_1503_ ;
wire \myexu/_1504_ ;
wire \myexu/_1505_ ;
wire \myexu/_1506_ ;
wire \myexu/_1507_ ;
wire \myexu/_1508_ ;
wire \myexu/_1509_ ;
wire \myexu/_1510_ ;
wire \myexu/_1511_ ;
wire \myexu/_1512_ ;
wire \myexu/_1513_ ;
wire \myexu/_1514_ ;
wire \myexu/_1515_ ;
wire \myexu/_1516_ ;
wire \myexu/_1517_ ;
wire \myexu/_1518_ ;
wire \myexu/_1519_ ;
wire \myexu/_1520_ ;
wire \myexu/_1521_ ;
wire \myexu/_1522_ ;
wire \myexu/_1523_ ;
wire \myexu/_1524_ ;
wire \myexu/_1525_ ;
wire \myexu/_1526_ ;
wire \myexu/_1527_ ;
wire \myexu/_1528_ ;
wire \myexu/_1529_ ;
wire \myexu/_1530_ ;
wire \myexu/_1531_ ;
wire \myexu/_1532_ ;
wire \myexu/_1533_ ;
wire \myexu/_1534_ ;
wire \myexu/_1535_ ;
wire \myexu/_1536_ ;
wire \myexu/_1537_ ;
wire \myexu/_1538_ ;
wire \myexu/_1539_ ;
wire \myexu/_1540_ ;
wire \myexu/_1541_ ;
wire \myexu/_1542_ ;
wire \myexu/_1543_ ;
wire \myexu/_1544_ ;
wire \myexu/_1545_ ;
wire \myexu/_1546_ ;
wire \myexu/_1547_ ;
wire \myexu/_1548_ ;
wire \myexu/_1549_ ;
wire \myexu/_1550_ ;
wire \myexu/_1551_ ;
wire \myexu/_1552_ ;
wire \myexu/_1553_ ;
wire \myexu/_1554_ ;
wire \myexu/_1555_ ;
wire \myexu/_1556_ ;
wire \myexu/_1557_ ;
wire \myexu/_1558_ ;
wire \myexu/_1559_ ;
wire \myexu/_1560_ ;
wire \myexu/_1561_ ;
wire \myexu/_1562_ ;
wire \myexu/_1563_ ;
wire \myexu/_1564_ ;
wire \myexu/_1565_ ;
wire \myexu/_1566_ ;
wire \myexu/_1567_ ;
wire \myexu/_1568_ ;
wire \myexu/_1569_ ;
wire \myexu/_1570_ ;
wire \myexu/_1571_ ;
wire \myexu/_1572_ ;
wire \myexu/_1573_ ;
wire \myexu/_1574_ ;
wire \myexu/_1575_ ;
wire \myexu/_1576_ ;
wire \myexu/_1577_ ;
wire \myexu/_1578_ ;
wire \myexu/_1579_ ;
wire \myexu/_1580_ ;
wire \myexu/_1581_ ;
wire \myexu/_1582_ ;
wire \myexu/_1583_ ;
wire \myexu/_1584_ ;
wire \myexu/_1585_ ;
wire \myexu/_1586_ ;
wire \myexu/_1587_ ;
wire \myexu/_1588_ ;
wire \myexu/_1589_ ;
wire \myexu/_1590_ ;
wire \myexu/_1591_ ;
wire \myexu/_1592_ ;
wire \myexu/_1593_ ;
wire \myexu/_1594_ ;
wire \myexu/_1595_ ;
wire \myexu/_1596_ ;
wire \myexu/_1597_ ;
wire \myexu/_1598_ ;
wire \myexu/_1599_ ;
wire \myexu/_1600_ ;
wire \myexu/_1601_ ;
wire \myexu/_1602_ ;
wire \myexu/_1603_ ;
wire \myexu/_1604_ ;
wire \myexu/_1605_ ;
wire \myexu/_1606_ ;
wire \myexu/_1607_ ;
wire \myexu/_1608_ ;
wire \myexu/_1609_ ;
wire \myexu/_1610_ ;
wire \myexu/_1611_ ;
wire \myexu/_1612_ ;
wire \myexu/_1613_ ;
wire \myexu/_1614_ ;
wire \myexu/_1615_ ;
wire \myexu/_1616_ ;
wire \myexu/_1617_ ;
wire \myexu/_1618_ ;
wire \myexu/_1619_ ;
wire \myexu/_1620_ ;
wire \myexu/_1621_ ;
wire \myexu/_1622_ ;
wire \myexu/_1623_ ;
wire \myexu/_1624_ ;
wire \myexu/_1625_ ;
wire \myexu/_1626_ ;
wire \myexu/_1627_ ;
wire \myexu/_1628_ ;
wire \myexu/_1629_ ;
wire \myexu/_1630_ ;
wire \myexu/_1631_ ;
wire \myexu/_1632_ ;
wire \myexu/_1633_ ;
wire \myexu/_1634_ ;
wire \myexu/_1635_ ;
wire \myexu/_1636_ ;
wire \myexu/_1637_ ;
wire \myexu/_1638_ ;
wire \myexu/_1639_ ;
wire \myexu/_1640_ ;
wire \myexu/_1641_ ;
wire \myexu/_1642_ ;
wire \myexu/_1643_ ;
wire \myexu/_1644_ ;
wire \myexu/_1645_ ;
wire \myexu/_1646_ ;
wire \myexu/_1647_ ;
wire \myexu/_1648_ ;
wire \myexu/_1649_ ;
wire \myexu/_1650_ ;
wire \myexu/_1651_ ;
wire \myexu/_1652_ ;
wire \myexu/_1653_ ;
wire \myexu/_1654_ ;
wire \myexu/_1655_ ;
wire \myexu/_1656_ ;
wire \myexu/_1657_ ;
wire \myexu/_1658_ ;
wire \myexu/_1659_ ;
wire \myexu/_1660_ ;
wire \myexu/_1661_ ;
wire \myexu/_1662_ ;
wire \myexu/_1663_ ;
wire \myexu/_1664_ ;
wire \myexu/_1665_ ;
wire \myexu/_1666_ ;
wire \myexu/_1667_ ;
wire \myexu/_1668_ ;
wire \myexu/_1669_ ;
wire \myexu/_1670_ ;
wire \myexu/_1671_ ;
wire \myexu/_1672_ ;
wire \myexu/_1673_ ;
wire \myexu/_1674_ ;
wire \myexu/_1675_ ;
wire \myexu/_1676_ ;
wire \myexu/_1677_ ;
wire \myexu/_1678_ ;
wire \myexu/_1679_ ;
wire \myexu/_1680_ ;
wire \myexu/_1681_ ;
wire \myexu/_1682_ ;
wire \myexu/_1683_ ;
wire \myexu/_1684_ ;
wire \myexu/_1685_ ;
wire \myexu/_1686_ ;
wire \myexu/_1687_ ;
wire \myexu/_1688_ ;
wire \myexu/_1689_ ;
wire \myexu/_1690_ ;
wire \myexu/_1691_ ;
wire \myexu/_1692_ ;
wire \myexu/_1693_ ;
wire \myexu/_1694_ ;
wire \myexu/_1695_ ;
wire \myexu/_1696_ ;
wire \myexu/_1697_ ;
wire \myexu/_1698_ ;
wire \myexu/_1699_ ;
wire \myexu/_1700_ ;
wire \myexu/_1701_ ;
wire \myexu/_1702_ ;
wire \myexu/_1703_ ;
wire \myexu/_1704_ ;
wire \myexu/_1705_ ;
wire \myexu/_1706_ ;
wire \myexu/_1707_ ;
wire \myexu/_1708_ ;
wire \myexu/_1709_ ;
wire \myexu/_1710_ ;
wire \myexu/_1711_ ;
wire \myexu/_1712_ ;
wire \myexu/_1713_ ;
wire \myexu/_1714_ ;
wire \myexu/_1715_ ;
wire \myexu/_1716_ ;
wire \myexu/_1717_ ;
wire \myexu/_1718_ ;
wire \myexu/_1719_ ;
wire \myexu/_1720_ ;
wire \myexu/_1721_ ;
wire \myexu/_1722_ ;
wire \myexu/_1723_ ;
wire \myexu/_1724_ ;
wire \myexu/_1725_ ;
wire \myexu/_1726_ ;
wire \myexu/_1727_ ;
wire \myexu/_1728_ ;
wire \myexu/_1729_ ;
wire \myexu/_1730_ ;
wire \myexu/_1731_ ;
wire \myexu/_1732_ ;
wire \myexu/_1733_ ;
wire \myexu/_1734_ ;
wire \myexu/_1735_ ;
wire \myexu/_1736_ ;
wire \myexu/_1737_ ;
wire \myexu/_1738_ ;
wire \myexu/_1739_ ;
wire \myexu/_1740_ ;
wire \myexu/_1741_ ;
wire \myexu/_1742_ ;
wire \myexu/_1743_ ;
wire \myexu/_1744_ ;
wire \myexu/_1745_ ;
wire \myexu/_1746_ ;
wire \myexu/_1747_ ;
wire \myexu/_1748_ ;
wire \myexu/_1749_ ;
wire \myexu/_1750_ ;
wire \myexu/_1751_ ;
wire \myexu/_1752_ ;
wire \myexu/_1753_ ;
wire \myexu/_1754_ ;
wire \myexu/_1755_ ;
wire \myexu/_1756_ ;
wire \myexu/_1757_ ;
wire \myexu/_1758_ ;
wire \myexu/_1759_ ;
wire \myexu/_1760_ ;
wire \myexu/_1761_ ;
wire \myexu/_1762_ ;
wire \myexu/_1763_ ;
wire \myexu/_1764_ ;
wire \myexu/_1765_ ;
wire \myexu/_1766_ ;
wire \myexu/_1767_ ;
wire \myexu/_1768_ ;
wire \myexu/_1769_ ;
wire \myexu/_1770_ ;
wire \myexu/_1771_ ;
wire \myexu/_1772_ ;
wire \myexu/_1773_ ;
wire \myexu/_1774_ ;
wire \myexu/_1775_ ;
wire \myexu/_1776_ ;
wire \myexu/_1777_ ;
wire \myexu/_1778_ ;
wire \myexu/_1779_ ;
wire \myexu/_1780_ ;
wire \myexu/_1781_ ;
wire \myexu/_1782_ ;
wire \myexu/_1783_ ;
wire \myexu/_1784_ ;
wire \myexu/_1785_ ;
wire \myexu/_1786_ ;
wire \myexu/_1787_ ;
wire \myexu/_1788_ ;
wire \myexu/_1789_ ;
wire \myexu/_1790_ ;
wire \myexu/_1791_ ;
wire \myexu/_1792_ ;
wire \myexu/_1793_ ;
wire \myexu/_1794_ ;
wire \myexu/_1795_ ;
wire \myexu/_1796_ ;
wire \myexu/_1797_ ;
wire \myexu/_1798_ ;
wire \myexu/_1799_ ;
wire \myexu/_1800_ ;
wire \myexu/_1801_ ;
wire \myexu/_1802_ ;
wire \myexu/_1803_ ;
wire \myexu/_1804_ ;
wire \myexu/_1805_ ;
wire \myexu/_1806_ ;
wire \myexu/_1807_ ;
wire \myexu/_1808_ ;
wire \myexu/_1809_ ;
wire \myexu/_1810_ ;
wire \myexu/_1811_ ;
wire \myexu/_1812_ ;
wire \myexu/_1813_ ;
wire \myexu/_1814_ ;
wire \myexu/_1815_ ;
wire \myexu/_1816_ ;
wire \myexu/_1817_ ;
wire \myexu/_1818_ ;
wire \myexu/_1819_ ;
wire \myexu/_1820_ ;
wire \myexu/_1821_ ;
wire \myexu/_1822_ ;
wire \myexu/_1823_ ;
wire \myexu/_1824_ ;
wire \myexu/_1825_ ;
wire \myexu/_1826_ ;
wire \myexu/_1827_ ;
wire \myexu/_1828_ ;
wire \myexu/_1829_ ;
wire \myexu/_1830_ ;
wire \myexu/_1831_ ;
wire \myexu/_1832_ ;
wire \myexu/_1833_ ;
wire \myexu/_1834_ ;
wire \myexu/_1835_ ;
wire \myexu/_1836_ ;
wire \myexu/_1837_ ;
wire \myexu/_1838_ ;
wire \myexu/_1839_ ;
wire \myexu/_1840_ ;
wire \myexu/_1841_ ;
wire \myexu/_1842_ ;
wire \myexu/_1843_ ;
wire \myexu/_1844_ ;
wire \myexu/_1845_ ;
wire \myexu/_1846_ ;
wire \myexu/_1847_ ;
wire \myexu/_1848_ ;
wire \myexu/_1849_ ;
wire \myexu/_1850_ ;
wire \myexu/_1851_ ;
wire \myexu/_1852_ ;
wire \myexu/_1853_ ;
wire \myexu/_1854_ ;
wire \myexu/_1855_ ;
wire \myexu/_1856_ ;
wire \myexu/_1857_ ;
wire \myexu/_1858_ ;
wire \myexu/_1859_ ;
wire \myexu/_1860_ ;
wire \myexu/_1861_ ;
wire \myexu/_1862_ ;
wire \myexu/_1863_ ;
wire \myexu/_1864_ ;
wire \myexu/_1865_ ;
wire \myexu/_1866_ ;
wire \myexu/_1867_ ;
wire \myexu/_1868_ ;
wire \myexu/_1869_ ;
wire \myexu/_1870_ ;
wire \myexu/_1871_ ;
wire \myexu/_1872_ ;
wire \myexu/_1873_ ;
wire \myexu/_1874_ ;
wire \myexu/_1875_ ;
wire \myexu/_1876_ ;
wire \myexu/_1877_ ;
wire \myexu/_1878_ ;
wire \myexu/_1879_ ;
wire \myexu/_1880_ ;
wire \myexu/_1881_ ;
wire \myexu/_1882_ ;
wire \myexu/_1883_ ;
wire \myexu/_1884_ ;
wire \myexu/_1885_ ;
wire \myexu/_1886_ ;
wire \myexu/_1887_ ;
wire \myexu/_1888_ ;
wire \myexu/_1889_ ;
wire \myexu/_1890_ ;
wire \myexu/_1891_ ;
wire \myexu/_1892_ ;
wire \myexu/_1893_ ;
wire \myexu/_1894_ ;
wire \myexu/_1895_ ;
wire \myexu/_1896_ ;
wire \myexu/_1897_ ;
wire \myexu/_1898_ ;
wire \myexu/_1899_ ;
wire \myexu/_1900_ ;
wire \myexu/_1901_ ;
wire \myexu/_1902_ ;
wire \myexu/_1903_ ;
wire \myexu/_1904_ ;
wire \myexu/_1905_ ;
wire \myexu/_1906_ ;
wire \myexu/_1907_ ;
wire \myexu/_1908_ ;
wire \myexu/_1909_ ;
wire \myexu/_1910_ ;
wire \myexu/_1911_ ;
wire \myexu/_1912_ ;
wire \myexu/_1913_ ;
wire \myexu/_1914_ ;
wire \myexu/_1915_ ;
wire \myexu/_1916_ ;
wire \myexu/_1917_ ;
wire \myexu/_1918_ ;
wire \myexu/_1919_ ;
wire \myexu/_1920_ ;
wire \myexu/_1921_ ;
wire \myexu/_1922_ ;
wire \myexu/_1923_ ;
wire \myexu/_1924_ ;
wire \myexu/_1925_ ;
wire \myexu/_1926_ ;
wire \myexu/_1927_ ;
wire \myexu/_1928_ ;
wire \myexu/_1929_ ;
wire \myexu/_1930_ ;
wire \myexu/_1931_ ;
wire \myexu/_1932_ ;
wire \myexu/_1933_ ;
wire \myexu/_1934_ ;
wire \myexu/_1935_ ;
wire \myexu/_1936_ ;
wire \myexu/_1937_ ;
wire \myexu/_1938_ ;
wire \myexu/_1939_ ;
wire \myexu/_1940_ ;
wire \myexu/_1941_ ;
wire \myexu/_1942_ ;
wire \myexu/_1943_ ;
wire \myexu/_1944_ ;
wire \myexu/_1945_ ;
wire \myexu/_1946_ ;
wire \myexu/_1947_ ;
wire \myexu/_1948_ ;
wire \myexu/_1949_ ;
wire \myexu/_1950_ ;
wire \myexu/_1951_ ;
wire \myexu/_1952_ ;
wire \myexu/_1953_ ;
wire \myexu/_1954_ ;
wire \myexu/_1955_ ;
wire \myexu/_1956_ ;
wire \myexu/_1957_ ;
wire \myexu/_1958_ ;
wire \myexu/_1959_ ;
wire \myexu/_1960_ ;
wire \myexu/_1961_ ;
wire \myexu/_1962_ ;
wire \myexu/_1963_ ;
wire \myexu/_1964_ ;
wire \myexu/_1965_ ;
wire \myexu/_1966_ ;
wire \myexu/_1967_ ;
wire \myexu/_1968_ ;
wire \myexu/_1969_ ;
wire \myexu/_1970_ ;
wire \myexu/_1971_ ;
wire \myexu/_1972_ ;
wire \myexu/_1973_ ;
wire \myexu/_1974_ ;
wire \myexu/_1975_ ;
wire \myexu/_1976_ ;
wire \myexu/_1977_ ;
wire \myexu/_1978_ ;
wire \myexu/_1979_ ;
wire \myexu/_1980_ ;
wire \myexu/_1981_ ;
wire \myexu/_1982_ ;
wire \myexu/_1983_ ;
wire \myexu/_1984_ ;
wire \myexu/_1985_ ;
wire \myexu/_1986_ ;
wire \myexu/_1987_ ;
wire \myexu/_1988_ ;
wire \myexu/_1989_ ;
wire \myexu/_1990_ ;
wire \myexu/_1991_ ;
wire \myexu/_1992_ ;
wire \myexu/_1993_ ;
wire \myexu/_1994_ ;
wire \myexu/_1995_ ;
wire \myexu/_1996_ ;
wire \myexu/_1997_ ;
wire \myexu/_1998_ ;
wire \myexu/_1999_ ;
wire \myexu/_2000_ ;
wire \myexu/_2001_ ;
wire \myexu/_2002_ ;
wire \myexu/_2003_ ;
wire \myexu/_2004_ ;
wire \myexu/_2005_ ;
wire \myexu/_2006_ ;
wire \myexu/_2007_ ;
wire \myexu/_2008_ ;
wire \myexu/_2009_ ;
wire \myexu/_2010_ ;
wire \myexu/_2011_ ;
wire \myexu/_2012_ ;
wire \myexu/_2013_ ;
wire \myexu/_2014_ ;
wire \myexu/_2015_ ;
wire \myexu/_2016_ ;
wire \myexu/_2017_ ;
wire \myexu/_2018_ ;
wire \myexu/_2019_ ;
wire \myexu/_2020_ ;
wire \myexu/_2021_ ;
wire \myexu/_2022_ ;
wire \myexu/_2023_ ;
wire \myexu/_2024_ ;
wire \myexu/_2025_ ;
wire \myexu/_2026_ ;
wire \myexu/_2027_ ;
wire \myexu/_2028_ ;
wire \myexu/_2029_ ;
wire \myexu/_2030_ ;
wire \myexu/_2031_ ;
wire \myexu/_2032_ ;
wire \myexu/_2033_ ;
wire \myexu/_2034_ ;
wire \myexu/_2035_ ;
wire \myexu/_2036_ ;
wire \myexu/_2037_ ;
wire \myexu/_2038_ ;
wire \myexu/_2039_ ;
wire \myexu/_2040_ ;
wire \myexu/_2041_ ;
wire \myexu/_2042_ ;
wire \myexu/_2043_ ;
wire \myexu/_2044_ ;
wire \myexu/_2045_ ;
wire \myexu/_2046_ ;
wire \myexu/_2047_ ;
wire \myexu/_2048_ ;
wire \myexu/_2049_ ;
wire \myexu/_2050_ ;
wire \myexu/_2051_ ;
wire \myexu/_2052_ ;
wire \myexu/_2053_ ;
wire \myexu/_2054_ ;
wire \myexu/_2055_ ;
wire \myexu/_2056_ ;
wire \myexu/_2057_ ;
wire \myexu/_2058_ ;
wire \myexu/_2059_ ;
wire \myexu/_2060_ ;
wire \myexu/_2061_ ;
wire \myexu/_2062_ ;
wire \myexu/_2063_ ;
wire \myexu/_2064_ ;
wire \myexu/_2065_ ;
wire \myexu/_2066_ ;
wire \myexu/_2067_ ;
wire \myexu/_2068_ ;
wire \myexu/_2069_ ;
wire \myexu/_2070_ ;
wire \myexu/_2071_ ;
wire \myexu/_2072_ ;
wire \myexu/_2073_ ;
wire \myexu/_2074_ ;
wire \myexu/_2075_ ;
wire \myexu/_2076_ ;
wire \myexu/_2077_ ;
wire \myexu/_2078_ ;
wire \myexu/_2079_ ;
wire \myexu/_2080_ ;
wire \myexu/_2081_ ;
wire \myexu/_2082_ ;
wire \myexu/_2083_ ;
wire \myexu/_2084_ ;
wire \myexu/_2085_ ;
wire \myexu/_2086_ ;
wire \myexu/_2087_ ;
wire \myexu/_2088_ ;
wire \myexu/_2089_ ;
wire \myexu/_2090_ ;
wire \myexu/_2091_ ;
wire \myexu/_2092_ ;
wire \myexu/_2093_ ;
wire \myexu/_2094_ ;
wire \myexu/_2095_ ;
wire \myexu/_2096_ ;
wire \myexu/_2097_ ;
wire \myexu/_2098_ ;
wire \myexu/_2099_ ;
wire \myexu/_2100_ ;
wire \myexu/_2101_ ;
wire \myexu/_2102_ ;
wire \myexu/_2103_ ;
wire \myexu/_2104_ ;
wire \myexu/_2105_ ;
wire \myexu/_2106_ ;
wire \myexu/_2107_ ;
wire \myexu/_2108_ ;
wire \myexu/_2109_ ;
wire \myexu/_2110_ ;
wire \myexu/_2111_ ;
wire \myexu/_2112_ ;
wire \myexu/_2113_ ;
wire \myexu/_2114_ ;
wire \myexu/_2115_ ;
wire \myexu/_2116_ ;
wire \myexu/_2117_ ;
wire \myexu/_2118_ ;
wire \myexu/_2119_ ;
wire \myexu/_2120_ ;
wire \myexu/_2121_ ;
wire \myexu/_2122_ ;
wire \myexu/_2123_ ;
wire \myexu/_2124_ ;
wire \myexu/_2125_ ;
wire \myexu/_2126_ ;
wire \myexu/_2127_ ;
wire \myexu/_2128_ ;
wire \myexu/_2129_ ;
wire \myexu/_2130_ ;
wire \myexu/_2131_ ;
wire \myexu/_2132_ ;
wire \myexu/_2133_ ;
wire \myexu/_2134_ ;
wire \myexu/_2135_ ;
wire \myexu/_2136_ ;
wire \myexu/_2137_ ;
wire \myexu/_2138_ ;
wire \myexu/_2139_ ;
wire \myexu/_2140_ ;
wire \myexu/_2141_ ;
wire \myexu/_2142_ ;
wire \myexu/_2143_ ;
wire \myexu/_2144_ ;
wire \myexu/_2145_ ;
wire \myexu/_2146_ ;
wire \myexu/_2147_ ;
wire \myexu/_2148_ ;
wire \myexu/_2149_ ;
wire \myexu/_2150_ ;
wire \myexu/_2151_ ;
wire \myexu/_2152_ ;
wire \myexu/_2153_ ;
wire \myexu/_2154_ ;
wire \myexu/_2155_ ;
wire \myexu/_2156_ ;
wire \myexu/_2157_ ;
wire \myexu/_2158_ ;
wire \myexu/_2159_ ;
wire \myexu/_2160_ ;
wire \myexu/_2161_ ;
wire \myexu/_2162_ ;
wire \myexu/_2163_ ;
wire \myexu/_2164_ ;
wire \myexu/_2165_ ;
wire \myexu/_2166_ ;
wire \myexu/_2167_ ;
wire \myexu/_2168_ ;
wire \myexu/_2169_ ;
wire \myexu/_2170_ ;
wire \myexu/_2171_ ;
wire \myexu/_2172_ ;
wire \myexu/_2173_ ;
wire \myexu/_2174_ ;
wire \myexu/_2175_ ;
wire \myexu/_2176_ ;
wire \myexu/_2177_ ;
wire \myexu/_2178_ ;
wire \myexu/_2179_ ;
wire \myexu/_2180_ ;
wire \myexu/_2181_ ;
wire \myexu/_2182_ ;
wire \myexu/_2183_ ;
wire \myexu/_2184_ ;
wire \myexu/_2185_ ;
wire \myexu/_2186_ ;
wire \myexu/_2187_ ;
wire \myexu/_2188_ ;
wire \myexu/_2189_ ;
wire \myexu/_2190_ ;
wire \myexu/_2191_ ;
wire \myexu/_2192_ ;
wire \myexu/_2193_ ;
wire \myexu/_2194_ ;
wire \myexu/_2195_ ;
wire \myexu/_2196_ ;
wire \myexu/_2197_ ;
wire \myexu/_2198_ ;
wire \myexu/_2199_ ;
wire \myexu/_2200_ ;
wire \myexu/_2201_ ;
wire \myexu/_2202_ ;
wire \myexu/_2203_ ;
wire \myexu/_2204_ ;
wire \myexu/_2205_ ;
wire \myexu/_2206_ ;
wire \myexu/_2207_ ;
wire \myexu/_2208_ ;
wire \myexu/_2209_ ;
wire \myexu/_2210_ ;
wire \myexu/_2211_ ;
wire \myexu/_2212_ ;
wire \myexu/_2213_ ;
wire \myexu/_2214_ ;
wire \myexu/_2215_ ;
wire \myexu/_2216_ ;
wire \myexu/_2217_ ;
wire \myexu/_2218_ ;
wire \myexu/_2219_ ;
wire \myexu/_2220_ ;
wire \myexu/_2221_ ;
wire \myexu/_2222_ ;
wire \myexu/_2223_ ;
wire \myexu/_2224_ ;
wire \myexu/_2225_ ;
wire \myexu/_2226_ ;
wire \myexu/_2227_ ;
wire \myexu/_2228_ ;
wire \myexu/_2229_ ;
wire \myexu/_2230_ ;
wire \myexu/_2231_ ;
wire \myexu/_2232_ ;
wire \myexu/_2233_ ;
wire \myexu/_2234_ ;
wire \myexu/_2235_ ;
wire \myexu/_2236_ ;
wire \myexu/_2237_ ;
wire \myexu/_2238_ ;
wire \myexu/_2239_ ;
wire \myexu/_2240_ ;
wire \myexu/_2241_ ;
wire \myexu/_2242_ ;
wire \myexu/_2243_ ;
wire \myexu/_2244_ ;
wire \myexu/_2245_ ;
wire \myexu/_2246_ ;
wire \myexu/_2247_ ;
wire \myexu/_2248_ ;
wire \myexu/_2249_ ;
wire \myexu/_2250_ ;
wire \myexu/_2251_ ;
wire \myexu/_2252_ ;
wire \myexu/_2253_ ;
wire \myexu/_2254_ ;
wire \myexu/_2255_ ;
wire \myexu/_2256_ ;
wire \myexu/_2257_ ;
wire \myexu/_2258_ ;
wire \myexu/_2259_ ;
wire \myexu/_2260_ ;
wire \myexu/_2261_ ;
wire \myexu/_2262_ ;
wire \myexu/_2263_ ;
wire \myexu/_2264_ ;
wire \myexu/_2265_ ;
wire \myexu/_2266_ ;
wire \myexu/_2267_ ;
wire \myexu/_2268_ ;
wire \myexu/_2269_ ;
wire \myexu/_2270_ ;
wire \myexu/_2271_ ;
wire \myexu/_2272_ ;
wire \myexu/_2273_ ;
wire \myexu/_2274_ ;
wire \myexu/_2275_ ;
wire \myexu/_2276_ ;
wire \myexu/_2277_ ;
wire \myexu/_2278_ ;
wire \myexu/_2279_ ;
wire \myexu/_2280_ ;
wire \myexu/_2281_ ;
wire \myexu/_2282_ ;
wire \myexu/_2283_ ;
wire \myexu/_2284_ ;
wire \myexu/_2285_ ;
wire \myexu/_2286_ ;
wire \myexu/_2287_ ;
wire \myexu/_2288_ ;
wire \myexu/_2289_ ;
wire \myexu/_2290_ ;
wire \myexu/_2291_ ;
wire \myexu/_2292_ ;
wire \myexu/_2293_ ;
wire \myexu/_2294_ ;
wire \myexu/_2295_ ;
wire \myexu/_2296_ ;
wire \myexu/_2297_ ;
wire \myexu/_2298_ ;
wire \myexu/_2299_ ;
wire \myexu/_2300_ ;
wire \myexu/_2301_ ;
wire \myexu/_2302_ ;
wire \myexu/_2303_ ;
wire \myexu/_2304_ ;
wire \myexu/_2305_ ;
wire \myexu/_2306_ ;
wire \myexu/_2307_ ;
wire \myexu/_2308_ ;
wire \myexu/_2309_ ;
wire \myexu/_2310_ ;
wire \myexu/_2311_ ;
wire \myexu/_2312_ ;
wire \myexu/_2313_ ;
wire \myexu/_2314_ ;
wire \myexu/_2315_ ;
wire \myexu/_2316_ ;
wire \myexu/_2317_ ;
wire \myexu/_2318_ ;
wire \myexu/_2319_ ;
wire \myexu/_2320_ ;
wire \myexu/_2321_ ;
wire \myexu/_2322_ ;
wire \myexu/_2323_ ;
wire \myexu/_2324_ ;
wire \myexu/_2325_ ;
wire \myexu/_2326_ ;
wire \myexu/_2327_ ;
wire \myexu/_2328_ ;
wire \myexu/_2329_ ;
wire \myexu/_2330_ ;
wire \myexu/_2331_ ;
wire \myexu/_2332_ ;
wire \myexu/_2333_ ;
wire \myexu/_2334_ ;
wire \myexu/_2335_ ;
wire \myexu/_2336_ ;
wire \myexu/_2337_ ;
wire \myexu/_2338_ ;
wire \myexu/_2339_ ;
wire \myexu/_2340_ ;
wire \myexu/_2341_ ;
wire \myexu/_2342_ ;
wire \myexu/_2343_ ;
wire \myexu/_2344_ ;
wire \myexu/_2345_ ;
wire \myexu/_2346_ ;
wire \myexu/_2347_ ;
wire \myexu/_2348_ ;
wire \myexu/_2349_ ;
wire \myexu/_2350_ ;
wire \myexu/_2351_ ;
wire \myexu/_2352_ ;
wire \myexu/_2353_ ;
wire \myexu/_2354_ ;
wire \myexu/_2355_ ;
wire \myexu/_2356_ ;
wire \myexu/_2357_ ;
wire \myexu/_2358_ ;
wire \myexu/_2359_ ;
wire \myexu/_2360_ ;
wire \myexu/_2361_ ;
wire \myexu/_2362_ ;
wire \myexu/_2363_ ;
wire \myexu/_2364_ ;
wire \myexu/_2365_ ;
wire \myexu/_2366_ ;
wire \myexu/_2367_ ;
wire \myexu/_2368_ ;
wire \myexu/_2369_ ;
wire \myexu/_2370_ ;
wire \myexu/_2371_ ;
wire \myexu/_2372_ ;
wire \myexu/_2373_ ;
wire \myexu/_2374_ ;
wire \myexu/_2375_ ;
wire \myexu/_2376_ ;
wire \myexu/_2377_ ;
wire \myexu/_2378_ ;
wire \myexu/_2379_ ;
wire \myexu/_2380_ ;
wire \myexu/_2381_ ;
wire \myexu/_2382_ ;
wire \myexu/_2383_ ;
wire \myexu/_2384_ ;
wire \myexu/_2385_ ;
wire \myexu/_2386_ ;
wire \myexu/_2387_ ;
wire \myexu/_2388_ ;
wire \myexu/_2389_ ;
wire \myexu/_2390_ ;
wire \myexu/_2391_ ;
wire \myexu/_2392_ ;
wire \myexu/_2393_ ;
wire \myexu/_2394_ ;
wire \myexu/_2395_ ;
wire \myexu/_2396_ ;
wire \myexu/_2397_ ;
wire \myexu/_2398_ ;
wire \myexu/_2399_ ;
wire \myexu/_2400_ ;
wire \myexu/_2401_ ;
wire \myexu/_2402_ ;
wire \myexu/_2403_ ;
wire \myexu/_2404_ ;
wire \myexu/_2405_ ;
wire \myexu/_2406_ ;
wire \myexu/_2407_ ;
wire \myexu/_2408_ ;
wire \myexu/_2409_ ;
wire \myexu/_2410_ ;
wire \myexu/_2411_ ;
wire \myexu/_2412_ ;
wire \myexu/_2413_ ;
wire \myexu/_2414_ ;
wire \myexu/_2415_ ;
wire \myexu/_2416_ ;
wire \myexu/_2417_ ;
wire \myexu/_2418_ ;
wire \myexu/_2419_ ;
wire \myexu/_2420_ ;
wire \myexu/_2421_ ;
wire \myexu/_2422_ ;
wire \myexu/_2423_ ;
wire \myexu/_2424_ ;
wire \myexu/_2425_ ;
wire \myexu/_2426_ ;
wire \myexu/_2427_ ;
wire \myexu/_2428_ ;
wire \myexu/_2429_ ;
wire \myexu/_2430_ ;
wire \myexu/_2431_ ;
wire \myexu/_2432_ ;
wire \myexu/_2433_ ;
wire \myexu/_2434_ ;
wire \myexu/_2435_ ;
wire \myexu/_2436_ ;
wire \myexu/_2437_ ;
wire \myexu/_2438_ ;
wire \myexu/_2439_ ;
wire \myexu/_2440_ ;
wire \myexu/_2441_ ;
wire \myexu/_2442_ ;
wire \myexu/_2443_ ;
wire \myexu/_2444_ ;
wire \myexu/_2445_ ;
wire \myexu/_2446_ ;
wire \myexu/_2447_ ;
wire \myexu/_2448_ ;
wire \myexu/_2449_ ;
wire \myexu/_2450_ ;
wire \myexu/_2451_ ;
wire \myexu/_2452_ ;
wire \myexu/_2453_ ;
wire \myexu/_2454_ ;
wire \myexu/_2455_ ;
wire \myexu/_2456_ ;
wire \myexu/_2457_ ;
wire \myexu/_2458_ ;
wire \myexu/_2459_ ;
wire \myexu/_2460_ ;
wire \myexu/_2461_ ;
wire \myexu/_2462_ ;
wire \myexu/_2463_ ;
wire \myexu/_2464_ ;
wire \myexu/_2465_ ;
wire \myexu/_2466_ ;
wire \myexu/_2467_ ;
wire \myexu/_2468_ ;
wire \myexu/_2469_ ;
wire \myexu/_2470_ ;
wire \myexu/_2471_ ;
wire \myexu/_2472_ ;
wire \myexu/_2473_ ;
wire \myexu/_2474_ ;
wire \myexu/_2475_ ;
wire \myexu/_2476_ ;
wire \myexu/_2477_ ;
wire \myexu/_2478_ ;
wire \myexu/_2479_ ;
wire \myexu/_2480_ ;
wire \myexu/_2481_ ;
wire \myexu/_2482_ ;
wire \myexu/_2483_ ;
wire \myexu/_2484_ ;
wire \myexu/_2485_ ;
wire \myexu/_2486_ ;
wire \myexu/_2487_ ;
wire \myexu/_2488_ ;
wire \myexu/_2489_ ;
wire \myexu/_2490_ ;
wire \myexu/_2491_ ;
wire \myexu/_2492_ ;
wire \myexu/_2493_ ;
wire \myexu/_2494_ ;
wire \myexu/_2495_ ;
wire \myexu/_2496_ ;
wire \myexu/_2497_ ;
wire \myexu/_2498_ ;
wire \myexu/_2499_ ;
wire \myexu/_2500_ ;
wire \myexu/_2501_ ;
wire \myexu/_2502_ ;
wire \myexu/_2503_ ;
wire \myexu/_2504_ ;
wire \myexu/_2505_ ;
wire \myexu/_2506_ ;
wire \myexu/_2507_ ;
wire \myexu/_2508_ ;
wire \myexu/_2509_ ;
wire \myexu/_2510_ ;
wire \myexu/_2511_ ;
wire \myexu/_2512_ ;
wire \myexu/_2513_ ;
wire \myexu/_2514_ ;
wire \myexu/_2515_ ;
wire \myexu/_2516_ ;
wire \myexu/_2517_ ;
wire \myexu/_2518_ ;
wire \myexu/_2519_ ;
wire \myexu/_2520_ ;
wire \myexu/_2521_ ;
wire \myexu/_2522_ ;
wire \myexu/_2523_ ;
wire \myexu/_2524_ ;
wire \myexu/_2525_ ;
wire \myexu/_2526_ ;
wire \myexu/_2527_ ;
wire \myexu/_2528_ ;
wire \myexu/_2529_ ;
wire \myexu/_2530_ ;
wire \myexu/_2531_ ;
wire \myexu/_2532_ ;
wire \myexu/_2533_ ;
wire \myexu/_2534_ ;
wire \myexu/_2535_ ;
wire \myexu/_2536_ ;
wire \myexu/_2537_ ;
wire \myexu/_2538_ ;
wire \myexu/_2539_ ;
wire \myexu/_2540_ ;
wire \myexu/_2541_ ;
wire \myexu/_2542_ ;
wire \myexu/_2543_ ;
wire \myexu/_2544_ ;
wire \myexu/_2545_ ;
wire \myexu/_2546_ ;
wire \myexu/_2547_ ;
wire \myexu/_2548_ ;
wire \myexu/_2549_ ;
wire \myexu/_2550_ ;
wire \myexu/_2551_ ;
wire \myexu/_2552_ ;
wire \myexu/_2553_ ;
wire \myexu/_2554_ ;
wire \myexu/_2555_ ;
wire \myexu/_2556_ ;
wire \myexu/_2557_ ;
wire \myexu/_2558_ ;
wire \myexu/_2559_ ;
wire \myexu/_2560_ ;
wire \myexu/_2561_ ;
wire \myexu/_2562_ ;
wire \myexu/_2563_ ;
wire \myexu/_2564_ ;
wire \myexu/_2565_ ;
wire \myexu/_2566_ ;
wire \myexu/_2567_ ;
wire \myexu/_2568_ ;
wire \myexu/_2569_ ;
wire \myexu/_2570_ ;
wire \myexu/_2571_ ;
wire \myexu/_2572_ ;
wire \myexu/_2573_ ;
wire \myexu/_2574_ ;
wire \myexu/_2575_ ;
wire \myexu/_2576_ ;
wire \myexu/_2577_ ;
wire \myexu/_2578_ ;
wire \myexu/_2579_ ;
wire \myexu/_2580_ ;
wire \myexu/_2581_ ;
wire \myexu/_2582_ ;
wire \myexu/_2583_ ;
wire \myexu/_2584_ ;
wire \myexu/_2585_ ;
wire \myexu/_2586_ ;
wire \myexu/_2587_ ;
wire \myexu/_2588_ ;
wire \myexu/_2589_ ;
wire \myexu/_2590_ ;
wire \myexu/_2591_ ;
wire \myexu/_2592_ ;
wire \myexu/_2593_ ;
wire \myexu/_2594_ ;
wire \myexu/_2595_ ;
wire \myexu/_2596_ ;
wire \myexu/_2597_ ;
wire \myexu/_2598_ ;
wire \myexu/_2599_ ;
wire \myexu/_2600_ ;
wire \myexu/_2601_ ;
wire \myexu/_2602_ ;
wire \myexu/_2603_ ;
wire \myexu/_2604_ ;
wire \myexu/_2605_ ;
wire \myexu/_2606_ ;
wire \myexu/_2607_ ;
wire \myexu/_2608_ ;
wire \myexu/_2609_ ;
wire \myexu/_2610_ ;
wire \myexu/_2611_ ;
wire \myexu/_2612_ ;
wire \myexu/_2613_ ;
wire \myexu/_2614_ ;
wire \myexu/_2615_ ;
wire \myexu/_2616_ ;
wire \myexu/_2617_ ;
wire \myexu/_2618_ ;
wire \myexu/_2619_ ;
wire \myexu/_2620_ ;
wire \myexu/_2621_ ;
wire \myexu/_2622_ ;
wire \myexu/_2623_ ;
wire \myexu/_2624_ ;
wire \myexu/_2625_ ;
wire \myexu/_2626_ ;
wire \myexu/_2627_ ;
wire \myexu/_2628_ ;
wire \myexu/_2629_ ;
wire \myexu/_2630_ ;
wire \myexu/_2631_ ;
wire \myexu/_2632_ ;
wire \myexu/_2633_ ;
wire \myexu/_2634_ ;
wire \myexu/_2635_ ;
wire \myexu/_2636_ ;
wire \myexu/_2637_ ;
wire \myexu/_2638_ ;
wire \myexu/_2639_ ;
wire \myexu/_2640_ ;
wire \myexu/_2641_ ;
wire \myexu/_2642_ ;
wire \myexu/_2643_ ;
wire \myexu/_2644_ ;
wire \myexu/_2645_ ;
wire \myexu/_2646_ ;
wire \myexu/_2647_ ;
wire \myexu/_2648_ ;
wire \myexu/_2649_ ;
wire \myexu/_2650_ ;
wire \myexu/_2651_ ;
wire \myexu/_2652_ ;
wire \myexu/_2653_ ;
wire \myexu/_2654_ ;
wire \myexu/_2655_ ;
wire \myexu/_2656_ ;
wire \myexu/_2657_ ;
wire \myexu/_2658_ ;
wire \myexu/_2659_ ;
wire \myexu/_2660_ ;
wire \myexu/_2661_ ;
wire \myexu/_2662_ ;
wire \myexu/_2663_ ;
wire \myexu/_2664_ ;
wire \myexu/_2665_ ;
wire \myexu/_2666_ ;
wire \myexu/_2667_ ;
wire \myexu/_2668_ ;
wire \myexu/_2669_ ;
wire \myexu/_2670_ ;
wire \myexu/_2671_ ;
wire \myexu/_2672_ ;
wire \myexu/_2673_ ;
wire \myexu/_2674_ ;
wire \myexu/_2675_ ;
wire \myexu/_2676_ ;
wire \myexu/_2677_ ;
wire \myexu/_2678_ ;
wire \myexu/_2679_ ;
wire \myexu/_2680_ ;
wire \myexu/_2681_ ;
wire \myexu/_2682_ ;
wire \myexu/_2683_ ;
wire \myexu/_2684_ ;
wire \myexu/_2685_ ;
wire \myexu/_2686_ ;
wire \myexu/_2687_ ;
wire \myexu/_2688_ ;
wire \myexu/_2689_ ;
wire \myexu/_2690_ ;
wire \myexu/_2691_ ;
wire \myexu/_2692_ ;
wire \myexu/_2693_ ;
wire \myexu/_2694_ ;
wire \myexu/_2695_ ;
wire \myexu/_2696_ ;
wire \myexu/_2697_ ;
wire \myexu/_2698_ ;
wire \myexu/_2699_ ;
wire \myexu/_2700_ ;
wire \myexu/_2701_ ;
wire \myexu/_2702_ ;
wire \myexu/_2703_ ;
wire \myexu/_2704_ ;
wire \myexu/_2705_ ;
wire \myexu/_2706_ ;
wire \myexu/_2707_ ;
wire \myexu/_2708_ ;
wire \myexu/_2709_ ;
wire \myexu/_2710_ ;
wire \myexu/_2711_ ;
wire \myexu/_2712_ ;
wire \myexu/_2713_ ;
wire \myexu/_2714_ ;
wire \myexu/_2715_ ;
wire \myexu/_2716_ ;
wire \myexu/_2717_ ;
wire \myexu/_2718_ ;
wire \myexu/_2719_ ;
wire \myexu/_2720_ ;
wire \myexu/_2721_ ;
wire \myexu/_2722_ ;
wire \myexu/_2723_ ;
wire \myexu/_2724_ ;
wire \myexu/_2725_ ;
wire \myexu/_2726_ ;
wire \myexu/_2727_ ;
wire \myexu/_2728_ ;
wire \myexu/_2729_ ;
wire \myexu/_2730_ ;
wire \myexu/_2731_ ;
wire \myexu/_2732_ ;
wire \myexu/_2733_ ;
wire \myexu/_2734_ ;
wire \myexu/_2735_ ;
wire \myexu/_2736_ ;
wire \myexu/_2737_ ;
wire \myexu/_2738_ ;
wire \myexu/_2739_ ;
wire \myexu/_2740_ ;
wire \myexu/_2741_ ;
wire \myexu/_2742_ ;
wire \myexu/_2743_ ;
wire \myexu/_2744_ ;
wire \myexu/_2745_ ;
wire \myexu/_2746_ ;
wire \myexu/_2747_ ;
wire \myexu/_2748_ ;
wire \myexu/_2749_ ;
wire \myexu/_2750_ ;
wire \myexu/_2751_ ;
wire \myexu/_2752_ ;
wire \myexu/_2753_ ;
wire \myexu/_2754_ ;
wire \myexu/_2755_ ;
wire \myexu/_2756_ ;
wire \myexu/_2757_ ;
wire \myexu/_2758_ ;
wire \myexu/_2759_ ;
wire \myexu/_2760_ ;
wire \myexu/_2761_ ;
wire \myexu/_2762_ ;
wire \myexu/_2763_ ;
wire \myexu/_2764_ ;
wire \myexu/_2765_ ;
wire \myexu/_2766_ ;
wire \myexu/_2767_ ;
wire \myexu/_2768_ ;
wire \myexu/_2769_ ;
wire \myexu/_2770_ ;
wire \myexu/_2771_ ;
wire \myexu/_2772_ ;
wire \myexu/_2773_ ;
wire \myexu/_2774_ ;
wire \myexu/_2775_ ;
wire \myexu/_2776_ ;
wire \myexu/_2777_ ;
wire \myexu/_2778_ ;
wire \myexu/_2779_ ;
wire \myexu/_2780_ ;
wire \myexu/_2781_ ;
wire \myexu/_2782_ ;
wire \myexu/_2783_ ;
wire \myexu/_2784_ ;
wire \myexu/_2785_ ;
wire \myexu/_2786_ ;
wire \myexu/_2787_ ;
wire \myexu/_2788_ ;
wire \myexu/_2789_ ;
wire \myexu/_2790_ ;
wire \myexu/_2791_ ;
wire \myexu/_2792_ ;
wire \myexu/_2793_ ;
wire \myexu/_2794_ ;
wire \myexu/_2795_ ;
wire \myexu/_2796_ ;
wire \myexu/_2797_ ;
wire \myexu/_2798_ ;
wire \myexu/_2799_ ;
wire \myexu/_2800_ ;
wire \myexu/_2801_ ;
wire \myexu/_2802_ ;
wire \myexu/_2803_ ;
wire \myexu/_2804_ ;
wire \myexu/_2805_ ;
wire \myexu/_2806_ ;
wire \myexu/_2807_ ;
wire \myexu/_2808_ ;
wire \myexu/_2809_ ;
wire \myexu/_2810_ ;
wire \myexu/_2811_ ;
wire \myexu/_2812_ ;
wire \myexu/_2813_ ;
wire \myexu/_2814_ ;
wire \myexu/_2815_ ;
wire \myexu/_2816_ ;
wire \myexu/_2817_ ;
wire \myexu/_2818_ ;
wire \myexu/_2819_ ;
wire \myexu/_2820_ ;
wire \myexu/_2821_ ;
wire \myexu/_2822_ ;
wire \myexu/_2823_ ;
wire \myexu/_2824_ ;
wire \myexu/_2825_ ;
wire \myexu/_2826_ ;
wire \myexu/_2827_ ;
wire \myexu/_2828_ ;
wire \myexu/_2829_ ;
wire \myexu/_2830_ ;
wire \myexu/_2831_ ;
wire \myexu/_2832_ ;
wire \myexu/_2833_ ;
wire \myexu/_2834_ ;
wire \myexu/_2835_ ;
wire \myexu/_2836_ ;
wire \myexu/_2837_ ;
wire \myexu/_2838_ ;
wire \myexu/_2839_ ;
wire \myexu/_2840_ ;
wire \myexu/_2841_ ;
wire \myexu/_2842_ ;
wire \myexu/_2843_ ;
wire \myexu/_2844_ ;
wire \myexu/_2845_ ;
wire \myexu/_2846_ ;
wire \myexu/_2847_ ;
wire \myexu/_2848_ ;
wire \myexu/_2849_ ;
wire \myexu/_2850_ ;
wire \myexu/_2851_ ;
wire \myexu/_2852_ ;
wire \myexu/_2853_ ;
wire \myexu/_2854_ ;
wire \myexu/_2855_ ;
wire \myexu/_2856_ ;
wire \myexu/_2857_ ;
wire \myexu/_2858_ ;
wire \myexu/_2859_ ;
wire \myexu/_2860_ ;
wire \myexu/_2861_ ;
wire \myexu/_2862_ ;
wire \myexu/_2863_ ;
wire \myexu/_2864_ ;
wire \myexu/_2865_ ;
wire \myexu/_2866_ ;
wire \myexu/_2867_ ;
wire \myexu/_2868_ ;
wire \myexu/_2869_ ;
wire \myexu/_2870_ ;
wire \myexu/_2871_ ;
wire \myexu/_2872_ ;
wire \myexu/_2873_ ;
wire \myexu/_2874_ ;
wire \myexu/_2875_ ;
wire \myexu/_2876_ ;
wire \myexu/_2877_ ;
wire \myexu/_2878_ ;
wire \myexu/_2879_ ;
wire \myexu/_2880_ ;
wire \myexu/_2881_ ;
wire \myexu/_2882_ ;
wire \myexu/_2883_ ;
wire \myexu/_2884_ ;
wire \myexu/_2885_ ;
wire \myexu/_2886_ ;
wire \myexu/myalu/_0000_ ;
wire \myexu/myalu/_0001_ ;
wire \myexu/myalu/_0002_ ;
wire \myexu/myalu/_0003_ ;
wire \myexu/myalu/_0004_ ;
wire \myexu/myalu/_0005_ ;
wire \myexu/myalu/_0006_ ;
wire \myexu/myalu/_0007_ ;
wire \myexu/myalu/_0008_ ;
wire \myexu/myalu/_0009_ ;
wire \myexu/myalu/_0010_ ;
wire \myexu/myalu/_0011_ ;
wire \myexu/myalu/_0012_ ;
wire \myexu/myalu/_0013_ ;
wire \myexu/myalu/_0014_ ;
wire \myexu/myalu/_0015_ ;
wire \myexu/myalu/_0016_ ;
wire \myexu/myalu/_0017_ ;
wire \myexu/myalu/_0018_ ;
wire \myexu/myalu/_0019_ ;
wire \myexu/myalu/_0020_ ;
wire \myexu/myalu/_0021_ ;
wire \myexu/myalu/_0022_ ;
wire \myexu/myalu/_0023_ ;
wire \myexu/myalu/_0024_ ;
wire \myexu/myalu/_0025_ ;
wire \myexu/myalu/_0026_ ;
wire \myexu/myalu/_0027_ ;
wire \myexu/myalu/_0028_ ;
wire \myexu/myalu/_0029_ ;
wire \myexu/myalu/_0030_ ;
wire \myexu/myalu/_0031_ ;
wire \myexu/myalu/_0032_ ;
wire \myexu/myalu/_0033_ ;
wire \myexu/myalu/_0034_ ;
wire \myexu/myalu/_0035_ ;
wire \myexu/myalu/_0036_ ;
wire \myexu/myalu/_0037_ ;
wire \myexu/myalu/_0038_ ;
wire \myexu/myalu/_0039_ ;
wire \myexu/myalu/_0040_ ;
wire \myexu/myalu/_0041_ ;
wire \myexu/myalu/_0042_ ;
wire \myexu/myalu/_0043_ ;
wire \myexu/myalu/_0044_ ;
wire \myexu/myalu/_0045_ ;
wire \myexu/myalu/_0046_ ;
wire \myexu/myalu/_0047_ ;
wire \myexu/myalu/_0048_ ;
wire \myexu/myalu/_0049_ ;
wire \myexu/myalu/_0050_ ;
wire \myexu/myalu/_0051_ ;
wire \myexu/myalu/_0052_ ;
wire \myexu/myalu/_0053_ ;
wire \myexu/myalu/_0054_ ;
wire \myexu/myalu/_0055_ ;
wire \myexu/myalu/_0056_ ;
wire \myexu/myalu/_0057_ ;
wire \myexu/myalu/_0058_ ;
wire \myexu/myalu/_0059_ ;
wire \myexu/myalu/_0060_ ;
wire \myexu/myalu/_0061_ ;
wire \myexu/myalu/_0062_ ;
wire \myexu/myalu/_0063_ ;
wire \myexu/myalu/_0064_ ;
wire \myexu/myalu/_0065_ ;
wire \myexu/myalu/_0066_ ;
wire \myexu/myalu/_0067_ ;
wire \myexu/myalu/_0068_ ;
wire \myexu/myalu/_0069_ ;
wire \myexu/myalu/_0070_ ;
wire \myexu/myalu/_0071_ ;
wire \myexu/myalu/_0072_ ;
wire \myexu/myalu/_0073_ ;
wire \myexu/myalu/_0074_ ;
wire \myexu/myalu/_0075_ ;
wire \myexu/myalu/_0076_ ;
wire \myexu/myalu/_0077_ ;
wire \myexu/myalu/_0078_ ;
wire \myexu/myalu/_0079_ ;
wire \myexu/myalu/_0080_ ;
wire \myexu/myalu/_0081_ ;
wire \myexu/myalu/_0082_ ;
wire \myexu/myalu/_0083_ ;
wire \myexu/myalu/_0084_ ;
wire \myexu/myalu/_0085_ ;
wire \myexu/myalu/_0086_ ;
wire \myexu/myalu/_0087_ ;
wire \myexu/myalu/_0088_ ;
wire \myexu/myalu/_0089_ ;
wire \myexu/myalu/_0090_ ;
wire \myexu/myalu/_0091_ ;
wire \myexu/myalu/_0092_ ;
wire \myexu/myalu/_0093_ ;
wire \myexu/myalu/_0094_ ;
wire \myexu/myalu/_0095_ ;
wire \myexu/myalu/_0096_ ;
wire \myexu/myalu/_0097_ ;
wire \myexu/myalu/_0098_ ;
wire \myexu/myalu/_0099_ ;
wire \myexu/myalu/_0100_ ;
wire \myexu/myalu/_0101_ ;
wire \myexu/myalu/_0102_ ;
wire \myexu/myalu/_0103_ ;
wire \myexu/myalu/_0104_ ;
wire \myexu/myalu/_0105_ ;
wire \myexu/myalu/_0106_ ;
wire \myexu/myalu/_0107_ ;
wire \myexu/myalu/_0108_ ;
wire \myexu/myalu/_0109_ ;
wire \myexu/myalu/_0110_ ;
wire \myexu/myalu/_0111_ ;
wire \myexu/myalu/_0112_ ;
wire \myexu/myalu/_0113_ ;
wire \myexu/myalu/_0114_ ;
wire \myexu/myalu/_0115_ ;
wire \myexu/myalu/_0116_ ;
wire \myexu/myalu/_0117_ ;
wire \myexu/myalu/_0118_ ;
wire \myexu/myalu/_0119_ ;
wire \myexu/myalu/_0120_ ;
wire \myexu/myalu/_0121_ ;
wire \myexu/myalu/_0122_ ;
wire \myexu/myalu/_0123_ ;
wire \myexu/myalu/_0124_ ;
wire \myexu/myalu/_0125_ ;
wire \myexu/myalu/_0126_ ;
wire \myexu/myalu/_0127_ ;
wire \myexu/myalu/_0128_ ;
wire \myexu/myalu/_0129_ ;
wire \myexu/myalu/_0130_ ;
wire \myexu/myalu/_0131_ ;
wire \myexu/myalu/_0132_ ;
wire \myexu/myalu/_0133_ ;
wire \myexu/myalu/_0134_ ;
wire \myexu/myalu/_0135_ ;
wire \myexu/myalu/_0136_ ;
wire \myexu/myalu/_0137_ ;
wire \myexu/myalu/_0138_ ;
wire \myexu/myalu/_0139_ ;
wire \myexu/myalu/_0140_ ;
wire \myexu/myalu/_0141_ ;
wire \myexu/myalu/_0142_ ;
wire \myexu/myalu/_0143_ ;
wire \myexu/myalu/_0144_ ;
wire \myexu/myalu/_0145_ ;
wire \myexu/myalu/_0146_ ;
wire \myexu/myalu/_0147_ ;
wire \myexu/myalu/_0148_ ;
wire \myexu/myalu/_0149_ ;
wire \myexu/myalu/_0150_ ;
wire \myexu/myalu/_0151_ ;
wire \myexu/myalu/_0152_ ;
wire \myexu/myalu/_0153_ ;
wire \myexu/myalu/_0154_ ;
wire \myexu/myalu/_0155_ ;
wire \myexu/myalu/_0156_ ;
wire \myexu/myalu/_0157_ ;
wire \myexu/myalu/_0158_ ;
wire \myexu/myalu/_0159_ ;
wire \myexu/myalu/_0160_ ;
wire \myexu/myalu/_0161_ ;
wire \myexu/myalu/_0162_ ;
wire \myexu/myalu/_0163_ ;
wire \myexu/myalu/_0164_ ;
wire \myexu/myalu/_0165_ ;
wire \myexu/myalu/_0166_ ;
wire \myexu/myalu/_0167_ ;
wire \myexu/myalu/_0168_ ;
wire \myexu/myalu/_0169_ ;
wire \myexu/myalu/_0170_ ;
wire \myexu/myalu/_0171_ ;
wire \myexu/myalu/_0172_ ;
wire \myexu/myalu/_0173_ ;
wire \myexu/myalu/_0174_ ;
wire \myexu/myalu/_0175_ ;
wire \myexu/myalu/_0176_ ;
wire \myexu/myalu/_0177_ ;
wire \myexu/myalu/_0178_ ;
wire \myexu/myalu/_0179_ ;
wire \myexu/myalu/_0180_ ;
wire \myexu/myalu/_0181_ ;
wire \myexu/myalu/_0182_ ;
wire \myexu/myalu/_0183_ ;
wire \myexu/myalu/_0184_ ;
wire \myexu/myalu/_0185_ ;
wire \myexu/myalu/_0186_ ;
wire \myexu/myalu/_0187_ ;
wire \myexu/myalu/_0188_ ;
wire \myexu/myalu/_0189_ ;
wire \myexu/myalu/_0190_ ;
wire \myexu/myalu/_0191_ ;
wire \myexu/myalu/_0192_ ;
wire \myexu/myalu/_0193_ ;
wire \myexu/myalu/_0194_ ;
wire \myexu/myalu/_0195_ ;
wire \myexu/myalu/_0196_ ;
wire \myexu/myalu/_0197_ ;
wire \myexu/myalu/_0198_ ;
wire \myexu/myalu/_0199_ ;
wire \myexu/myalu/_0200_ ;
wire \myexu/myalu/_0201_ ;
wire \myexu/myalu/_0202_ ;
wire \myexu/myalu/_0203_ ;
wire \myexu/myalu/_0204_ ;
wire \myexu/myalu/_0205_ ;
wire \myexu/myalu/_0206_ ;
wire \myexu/myalu/_0207_ ;
wire \myexu/myalu/_0208_ ;
wire \myexu/myalu/_0209_ ;
wire \myexu/myalu/_0210_ ;
wire \myexu/myalu/_0211_ ;
wire \myexu/myalu/_0212_ ;
wire \myexu/myalu/_0213_ ;
wire \myexu/myalu/_0214_ ;
wire \myexu/myalu/_0215_ ;
wire \myexu/myalu/_0216_ ;
wire \myexu/myalu/_0217_ ;
wire \myexu/myalu/_0218_ ;
wire \myexu/myalu/_0219_ ;
wire \myexu/myalu/_0220_ ;
wire \myexu/myalu/_0221_ ;
wire \myexu/myalu/_0222_ ;
wire \myexu/myalu/_0223_ ;
wire \myexu/myalu/_0224_ ;
wire \myexu/myalu/_0225_ ;
wire \myexu/myalu/_0226_ ;
wire \myexu/myalu/_0227_ ;
wire \myexu/myalu/_0228_ ;
wire \myexu/myalu/_0229_ ;
wire \myexu/myalu/_0230_ ;
wire \myexu/myalu/_0231_ ;
wire \myexu/myalu/_0232_ ;
wire \myexu/myalu/_0233_ ;
wire \myexu/myalu/_0234_ ;
wire \myexu/myalu/_0235_ ;
wire \myexu/myalu/_0236_ ;
wire \myexu/myalu/_0237_ ;
wire \myexu/myalu/_0238_ ;
wire \myexu/myalu/_0239_ ;
wire \myexu/myalu/_0240_ ;
wire \myexu/myalu/_0241_ ;
wire \myexu/myalu/_0242_ ;
wire \myexu/myalu/_0243_ ;
wire \myexu/myalu/_0244_ ;
wire \myexu/myalu/_0245_ ;
wire \myexu/myalu/_0246_ ;
wire \myexu/myalu/_0247_ ;
wire \myexu/myalu/_0248_ ;
wire \myexu/myalu/_0249_ ;
wire \myexu/myalu/_0250_ ;
wire \myexu/myalu/_0251_ ;
wire \myexu/myalu/_0252_ ;
wire \myexu/myalu/_0253_ ;
wire \myexu/myalu/_0254_ ;
wire \myexu/myalu/_0255_ ;
wire \myexu/myalu/_0256_ ;
wire \myexu/myalu/_0257_ ;
wire \myexu/myalu/_0258_ ;
wire \myexu/myalu/_0259_ ;
wire \myexu/myalu/_0260_ ;
wire \myexu/myalu/_0261_ ;
wire \myexu/myalu/_0262_ ;
wire \myexu/myalu/_0263_ ;
wire \myexu/myalu/_0264_ ;
wire \myexu/myalu/_0265_ ;
wire \myexu/myalu/_0266_ ;
wire \myexu/myalu/_0267_ ;
wire \myexu/myalu/_0268_ ;
wire \myexu/myalu/_0269_ ;
wire \myexu/myalu/_0270_ ;
wire \myexu/myalu/_0271_ ;
wire \myexu/myalu/_0272_ ;
wire \myexu/myalu/_0273_ ;
wire \myexu/myalu/_0274_ ;
wire \myexu/myalu/_0275_ ;
wire \myexu/myalu/_0276_ ;
wire \myexu/myalu/_0277_ ;
wire \myexu/myalu/_0278_ ;
wire \myexu/myalu/_0279_ ;
wire \myexu/myalu/_0280_ ;
wire \myexu/myalu/_0281_ ;
wire \myexu/myalu/_0282_ ;
wire \myexu/myalu/_0283_ ;
wire \myexu/myalu/_0284_ ;
wire \myexu/myalu/_0285_ ;
wire \myexu/myalu/_0286_ ;
wire \myexu/myalu/_0287_ ;
wire \myexu/myalu/_0288_ ;
wire \myexu/myalu/_0289_ ;
wire \myexu/myalu/_0290_ ;
wire \myexu/myalu/_0291_ ;
wire \myexu/myalu/_0292_ ;
wire \myexu/myalu/_0293_ ;
wire \myexu/myalu/_0294_ ;
wire \myexu/myalu/_0295_ ;
wire \myexu/myalu/_0296_ ;
wire \myexu/myalu/_0297_ ;
wire \myexu/myalu/_0298_ ;
wire \myexu/myalu/_0299_ ;
wire \myexu/myalu/_0300_ ;
wire \myexu/myalu/_0301_ ;
wire \myexu/myalu/_0302_ ;
wire \myexu/myalu/_0303_ ;
wire \myexu/myalu/_0304_ ;
wire \myexu/myalu/_0305_ ;
wire \myexu/myalu/_0306_ ;
wire \myexu/myalu/_0307_ ;
wire \myexu/myalu/_0308_ ;
wire \myexu/myalu/_0309_ ;
wire \myexu/myalu/_0310_ ;
wire \myexu/myalu/_0311_ ;
wire \myexu/myalu/_0312_ ;
wire \myexu/myalu/_0313_ ;
wire \myexu/myalu/_0314_ ;
wire \myexu/myalu/_0315_ ;
wire \myexu/myalu/_0316_ ;
wire \myexu/myalu/_0317_ ;
wire \myexu/myalu/_0318_ ;
wire \myexu/myalu/_0319_ ;
wire \myexu/myalu/_0320_ ;
wire \myexu/myalu/_0321_ ;
wire \myexu/myalu/_0322_ ;
wire \myexu/myalu/_0323_ ;
wire \myexu/myalu/_0324_ ;
wire \myexu/myalu/_0325_ ;
wire \myexu/myalu/_0326_ ;
wire \myexu/myalu/_0327_ ;
wire \myexu/myalu/_0328_ ;
wire \myexu/myalu/_0329_ ;
wire \myexu/myalu/_0330_ ;
wire \myexu/myalu/_0331_ ;
wire \myexu/myalu/_0332_ ;
wire \myexu/myalu/_0333_ ;
wire \myexu/myalu/_0334_ ;
wire \myexu/myalu/_0335_ ;
wire \myexu/myalu/_0336_ ;
wire \myexu/myalu/_0337_ ;
wire \myexu/myalu/_0338_ ;
wire \myexu/myalu/_0339_ ;
wire \myexu/myalu/_0340_ ;
wire \myexu/myalu/_0341_ ;
wire \myexu/myalu/_0342_ ;
wire \myexu/myalu/_0343_ ;
wire \myexu/myalu/_0344_ ;
wire \myexu/myalu/_0345_ ;
wire \myexu/myalu/_0346_ ;
wire \myexu/myalu/_0347_ ;
wire \myexu/myalu/_0348_ ;
wire \myexu/myalu/_0349_ ;
wire \myexu/myalu/_0350_ ;
wire \myexu/myalu/_0351_ ;
wire \myexu/myalu/_0352_ ;
wire \myexu/myalu/_0353_ ;
wire \myexu/myalu/_0354_ ;
wire \myexu/myalu/_0355_ ;
wire \myexu/myalu/_0356_ ;
wire \myexu/myalu/_0357_ ;
wire \myexu/myalu/_0358_ ;
wire \myexu/myalu/_0359_ ;
wire \myexu/myalu/_0360_ ;
wire \myexu/myalu/_0361_ ;
wire \myexu/myalu/_0362_ ;
wire \myexu/myalu/_0363_ ;
wire \myexu/myalu/_0364_ ;
wire \myexu/myalu/_0365_ ;
wire \myexu/myalu/_0366_ ;
wire \myexu/myalu/_0367_ ;
wire \myexu/myalu/_0368_ ;
wire \myexu/myalu/_0369_ ;
wire \myexu/myalu/_0370_ ;
wire \myexu/myalu/_0371_ ;
wire \myexu/myalu/_0372_ ;
wire \myexu/myalu/_0373_ ;
wire \myexu/myalu/_0374_ ;
wire \myexu/myalu/_0375_ ;
wire \myexu/myalu/_0376_ ;
wire \myexu/myalu/_0377_ ;
wire \myexu/myalu/_0378_ ;
wire \myexu/myalu/_0379_ ;
wire \myexu/myalu/_0380_ ;
wire \myexu/myalu/_0381_ ;
wire \myexu/myalu/_0382_ ;
wire \myexu/myalu/_0383_ ;
wire \myexu/myalu/_0384_ ;
wire \myexu/myalu/_0385_ ;
wire \myexu/myalu/_0386_ ;
wire \myexu/myalu/_0387_ ;
wire \myexu/myalu/_0388_ ;
wire \myexu/myalu/_0389_ ;
wire \myexu/myalu/_0390_ ;
wire \myexu/myalu/_0391_ ;
wire \myexu/myalu/_0392_ ;
wire \myexu/myalu/_0393_ ;
wire \myexu/myalu/_0394_ ;
wire \myexu/myalu/_0395_ ;
wire \myexu/myalu/_0396_ ;
wire \myexu/myalu/_0397_ ;
wire \myexu/myalu/_0398_ ;
wire \myexu/myalu/_0399_ ;
wire \myexu/myalu/_0400_ ;
wire \myexu/myalu/_0401_ ;
wire \myexu/myalu/_0402_ ;
wire \myexu/myalu/_0403_ ;
wire \myexu/myalu/_0404_ ;
wire \myexu/myalu/_0405_ ;
wire \myexu/myalu/_0406_ ;
wire \myexu/myalu/_0407_ ;
wire \myexu/myalu/_0408_ ;
wire \myexu/myalu/_0409_ ;
wire \myexu/myalu/_0410_ ;
wire \myexu/myalu/_0411_ ;
wire \myexu/myalu/_0412_ ;
wire \myexu/myalu/_0413_ ;
wire \myexu/myalu/_0414_ ;
wire \myexu/myalu/_0415_ ;
wire \myexu/myalu/_0416_ ;
wire \myexu/myalu/_0417_ ;
wire \myexu/myalu/_0418_ ;
wire \myexu/myalu/_0419_ ;
wire \myexu/myalu/_0420_ ;
wire \myexu/myalu/_0421_ ;
wire \myexu/myalu/_0422_ ;
wire \myexu/myalu/_0423_ ;
wire \myexu/myalu/_0424_ ;
wire \myexu/myalu/_0425_ ;
wire \myexu/myalu/_0426_ ;
wire \myexu/myalu/_0427_ ;
wire \myexu/myalu/_0428_ ;
wire \myexu/myalu/_0429_ ;
wire \myexu/myalu/_0430_ ;
wire \myexu/myalu/_0431_ ;
wire \myexu/myalu/_0432_ ;
wire \myexu/myalu/_0433_ ;
wire \myexu/myalu/_0434_ ;
wire \myexu/myalu/_0435_ ;
wire \myexu/myalu/_0436_ ;
wire \myexu/myalu/_0437_ ;
wire \myexu/myalu/_0438_ ;
wire \myexu/myalu/_0439_ ;
wire \myexu/myalu/_0440_ ;
wire \myexu/myalu/_0441_ ;
wire \myexu/myalu/_0442_ ;
wire \myexu/myalu/_0443_ ;
wire \myexu/myalu/_0444_ ;
wire \myexu/myalu/_0445_ ;
wire \myexu/myalu/_0446_ ;
wire \myexu/myalu/_0447_ ;
wire \myexu/myalu/_0448_ ;
wire \myexu/myalu/_0449_ ;
wire \myexu/myalu/_0450_ ;
wire \myexu/myalu/_0451_ ;
wire \myexu/myalu/_0452_ ;
wire \myexu/myalu/_0453_ ;
wire \myexu/myalu/_0454_ ;
wire \myexu/myalu/_0455_ ;
wire \myexu/myalu/_0456_ ;
wire \myexu/myalu/_0457_ ;
wire \myexu/myalu/_0458_ ;
wire \myexu/myalu/_0459_ ;
wire \myexu/myalu/_0460_ ;
wire \myexu/myalu/_0461_ ;
wire \myexu/myalu/_0462_ ;
wire \myexu/myalu/_0463_ ;
wire \myexu/myalu/_0464_ ;
wire \myexu/myalu/_0465_ ;
wire \myexu/myalu/_0466_ ;
wire \myexu/myalu/_0467_ ;
wire \myexu/myalu/_0468_ ;
wire \myexu/myalu/_0469_ ;
wire \myexu/myalu/_0470_ ;
wire \myexu/myalu/_0471_ ;
wire \myexu/myalu/_0472_ ;
wire \myexu/myalu/_0473_ ;
wire \myexu/myalu/_0474_ ;
wire \myexu/myalu/_0475_ ;
wire \myexu/myalu/_0476_ ;
wire \myexu/myalu/_0477_ ;
wire \myexu/myalu/_0478_ ;
wire \myexu/myalu/_0479_ ;
wire \myexu/myalu/_0480_ ;
wire \myexu/myalu/_0481_ ;
wire \myexu/myalu/_0482_ ;
wire \myexu/myalu/_0483_ ;
wire \myexu/myalu/_0484_ ;
wire \myexu/myalu/_0485_ ;
wire \myexu/myalu/_0486_ ;
wire \myexu/myalu/_0487_ ;
wire \myexu/myalu/_0488_ ;
wire \myexu/myalu/_0489_ ;
wire \myexu/myalu/_0490_ ;
wire \myexu/myalu/_0491_ ;
wire \myexu/myalu/_0492_ ;
wire \myexu/myalu/_0493_ ;
wire \myexu/myalu/_0494_ ;
wire \myexu/myalu/_0495_ ;
wire \myexu/myalu/_0496_ ;
wire \myexu/myalu/_0497_ ;
wire \myexu/myalu/_0498_ ;
wire \myexu/myalu/_0499_ ;
wire \myexu/myalu/_0500_ ;
wire \myexu/myalu/_0501_ ;
wire \myexu/myalu/_0502_ ;
wire \myexu/myalu/_0503_ ;
wire \myexu/myalu/_0504_ ;
wire \myexu/myalu/_0505_ ;
wire \myexu/myalu/_0506_ ;
wire \myexu/myalu/_0507_ ;
wire \myexu/myalu/_0508_ ;
wire \myexu/myalu/_0509_ ;
wire \myexu/myalu/_0510_ ;
wire \myexu/myalu/_0511_ ;
wire \myexu/myalu/_0512_ ;
wire \myexu/myalu/_0513_ ;
wire \myexu/myalu/_0514_ ;
wire \myexu/myalu/_0515_ ;
wire \myexu/myalu/_0516_ ;
wire \myexu/myalu/_0517_ ;
wire \myexu/myalu/_0518_ ;
wire \myexu/myalu/_0519_ ;
wire \myexu/myalu/_0520_ ;
wire \myexu/myalu/_0521_ ;
wire \myexu/myalu/_0522_ ;
wire \myexu/myalu/_0523_ ;
wire \myexu/myalu/_0524_ ;
wire \myexu/myalu/_0525_ ;
wire \myexu/myalu/_0526_ ;
wire \myexu/myalu/_0527_ ;
wire \myexu/myalu/_0528_ ;
wire \myexu/myalu/_0529_ ;
wire \myexu/myalu/_0530_ ;
wire \myexu/myalu/_0531_ ;
wire \myexu/myalu/_0532_ ;
wire \myexu/myalu/_0533_ ;
wire \myexu/myalu/_0534_ ;
wire \myexu/myalu/_0535_ ;
wire \myexu/myalu/_0536_ ;
wire \myexu/myalu/_0537_ ;
wire \myexu/myalu/_0538_ ;
wire \myexu/myalu/_0539_ ;
wire \myexu/myalu/_0540_ ;
wire \myexu/myalu/_0541_ ;
wire \myexu/myalu/_0542_ ;
wire \myexu/myalu/_0543_ ;
wire \myexu/myalu/_0544_ ;
wire \myexu/myalu/_0545_ ;
wire \myexu/myalu/_0546_ ;
wire \myexu/myalu/_0547_ ;
wire \myexu/myalu/_0548_ ;
wire \myexu/myalu/_0549_ ;
wire \myexu/myalu/_0550_ ;
wire \myexu/myalu/_0551_ ;
wire \myexu/myalu/_0552_ ;
wire \myexu/myalu/_0553_ ;
wire \myexu/myalu/_0554_ ;
wire \myexu/myalu/_0555_ ;
wire \myexu/myalu/_0556_ ;
wire \myexu/myalu/_0557_ ;
wire \myexu/myalu/_0558_ ;
wire \myexu/myalu/_0559_ ;
wire \myexu/myalu/_0560_ ;
wire \myexu/myalu/_0561_ ;
wire \myexu/myalu/_0562_ ;
wire \myexu/myalu/_0563_ ;
wire \myexu/myalu/_0564_ ;
wire \myexu/myalu/_0565_ ;
wire \myexu/myalu/_0566_ ;
wire \myexu/myalu/_0567_ ;
wire \myexu/myalu/_0568_ ;
wire \myexu/myalu/_0569_ ;
wire \myexu/myalu/_0570_ ;
wire \myexu/myalu/_0571_ ;
wire \myexu/myalu/_0572_ ;
wire \myexu/myalu/_0573_ ;
wire \myexu/myalu/_0574_ ;
wire \myexu/myalu/_0575_ ;
wire \myexu/myalu/_0576_ ;
wire \myexu/myalu/_0577_ ;
wire \myexu/myalu/_0578_ ;
wire \myexu/myalu/_0579_ ;
wire \myexu/myalu/_0580_ ;
wire \myexu/myalu/_0581_ ;
wire \myexu/myalu/_0582_ ;
wire \myexu/myalu/_0583_ ;
wire \myexu/myalu/_0584_ ;
wire \myexu/myalu/_0585_ ;
wire \myexu/myalu/_0586_ ;
wire \myexu/myalu/_0587_ ;
wire \myexu/myalu/_0588_ ;
wire \myexu/myalu/_0589_ ;
wire \myexu/myalu/_0590_ ;
wire \myexu/myalu/_0591_ ;
wire \myexu/myalu/_0592_ ;
wire \myexu/myalu/_0593_ ;
wire \myexu/myalu/_0594_ ;
wire \myexu/myalu/_0595_ ;
wire \myexu/myalu/_0596_ ;
wire \myexu/myalu/_0597_ ;
wire \myexu/myalu/_0598_ ;
wire \myexu/myalu/_0599_ ;
wire \myexu/myalu/_0600_ ;
wire \myexu/myalu/_0601_ ;
wire \myexu/myalu/_0602_ ;
wire \myexu/myalu/_0603_ ;
wire \myexu/myalu/_0604_ ;
wire \myexu/myalu/_0605_ ;
wire \myexu/myalu/_0606_ ;
wire \myexu/myalu/_0607_ ;
wire \myexu/myalu/_0608_ ;
wire \myexu/myalu/_0609_ ;
wire \myexu/myalu/_0610_ ;
wire \myexu/myalu/_0611_ ;
wire \myexu/myalu/_0612_ ;
wire \myexu/myalu/_0613_ ;
wire \myexu/myalu/_0614_ ;
wire \myexu/myalu/_0615_ ;
wire \myexu/myalu/_0616_ ;
wire \myexu/myalu/_0617_ ;
wire \myexu/myalu/_0618_ ;
wire \myexu/myalu/_0619_ ;
wire \myexu/myalu/_0620_ ;
wire \myexu/myalu/_0621_ ;
wire \myexu/myalu/_0622_ ;
wire \myexu/myalu/_0623_ ;
wire \myexu/myalu/_0624_ ;
wire \myexu/myalu/_0625_ ;
wire \myexu/myalu/_0626_ ;
wire \myexu/myalu/_0627_ ;
wire \myexu/myalu/_0628_ ;
wire \myexu/myalu/_0629_ ;
wire \myexu/myalu/_0630_ ;
wire \myexu/myalu/_0631_ ;
wire \myexu/myalu/_0632_ ;
wire \myexu/myalu/_0633_ ;
wire \myexu/myalu/_0634_ ;
wire \myexu/myalu/_0635_ ;
wire \myexu/myalu/_0636_ ;
wire \myexu/myalu/_0637_ ;
wire \myexu/myalu/_0638_ ;
wire \myexu/myalu/_0639_ ;
wire \myexu/myalu/_0640_ ;
wire \myexu/myalu/_0641_ ;
wire \myexu/myalu/_0642_ ;
wire \myexu/myalu/_0643_ ;
wire \myexu/myalu/_0644_ ;
wire \myexu/myalu/_0645_ ;
wire \myexu/myalu/_0646_ ;
wire \myexu/myalu/_0647_ ;
wire \myexu/myalu/_0648_ ;
wire \myexu/myalu/_0649_ ;
wire \myexu/myalu/_0650_ ;
wire \myexu/myalu/_0651_ ;
wire \myexu/myalu/_0652_ ;
wire \myexu/myalu/_0653_ ;
wire \myexu/myalu/_0654_ ;
wire \myexu/myalu/_0655_ ;
wire \myexu/myalu/_0656_ ;
wire \myexu/myalu/_0657_ ;
wire \myexu/myalu/_0658_ ;
wire \myexu/myalu/_0659_ ;
wire \myexu/myalu/_0660_ ;
wire \myexu/myalu/_0661_ ;
wire \myexu/myalu/_0662_ ;
wire \myexu/myalu/_0663_ ;
wire \myexu/myalu/_0664_ ;
wire \myexu/myalu/_0665_ ;
wire \myexu/myalu/_0666_ ;
wire \myexu/myalu/_0667_ ;
wire \myexu/myalu/_0668_ ;
wire \myexu/myalu/_0669_ ;
wire \myexu/myalu/_0670_ ;
wire \myexu/myalu/_0671_ ;
wire \myexu/myalu/_0672_ ;
wire \myexu/myalu/_0673_ ;
wire \myexu/myalu/_0674_ ;
wire \myexu/myalu/_0675_ ;
wire \myexu/myalu/_0676_ ;
wire \myexu/myalu/_0677_ ;
wire \myexu/myalu/_0678_ ;
wire \myexu/myalu/_0679_ ;
wire \myexu/myalu/_0680_ ;
wire \myexu/myalu/_0681_ ;
wire \myexu/myalu/_0682_ ;
wire \myexu/myalu/_0683_ ;
wire \myexu/myalu/_0684_ ;
wire \myexu/myalu/_0685_ ;
wire \myexu/myalu/_0686_ ;
wire \myexu/myalu/_0687_ ;
wire \myexu/myalu/_0688_ ;
wire \myexu/myalu/_0689_ ;
wire \myexu/myalu/_0690_ ;
wire \myexu/myalu/_0691_ ;
wire \myexu/myalu/_0692_ ;
wire \myexu/myalu/_0693_ ;
wire \myexu/myalu/_0694_ ;
wire \myexu/myalu/_0695_ ;
wire \myexu/myalu/_0696_ ;
wire \myexu/myalu/_0697_ ;
wire \myexu/myalu/_0698_ ;
wire \myexu/myalu/_0699_ ;
wire \myexu/myalu/_0700_ ;
wire \myexu/myalu/_0701_ ;
wire \myexu/myalu/_0702_ ;
wire \myexu/myalu/_0703_ ;
wire \myexu/myalu/_0704_ ;
wire \myexu/myalu/_0705_ ;
wire \myexu/myalu/_0706_ ;
wire \myexu/myalu/_0707_ ;
wire \myexu/myalu/_0708_ ;
wire \myexu/myalu/_0709_ ;
wire \myexu/myalu/_0710_ ;
wire \myexu/myalu/_0711_ ;
wire \myexu/myalu/_0712_ ;
wire \myexu/myalu/_0713_ ;
wire \myexu/myalu/_0714_ ;
wire \myexu/myalu/_0715_ ;
wire \myexu/myalu/_0716_ ;
wire \myexu/myalu/_0717_ ;
wire \myexu/myalu/_0718_ ;
wire \myexu/myalu/_0719_ ;
wire \myexu/myalu/_0720_ ;
wire \myexu/myalu/_0721_ ;
wire \myexu/myalu/_0722_ ;
wire \myexu/myalu/_0723_ ;
wire \myexu/myalu/_0724_ ;
wire \myexu/myalu/_0725_ ;
wire \myexu/myalu/_0726_ ;
wire \myexu/myalu/_0727_ ;
wire \myexu/myalu/_0728_ ;
wire \myexu/myalu/_0729_ ;
wire \myexu/myalu/_0730_ ;
wire \myexu/myalu/_0731_ ;
wire \myexu/myalu/_0732_ ;
wire \myexu/myalu/_0733_ ;
wire \myexu/myalu/_0734_ ;
wire \myexu/myalu/_0735_ ;
wire \myexu/myalu/_0736_ ;
wire \myexu/myalu/_0737_ ;
wire \myexu/myalu/_0738_ ;
wire \myexu/myalu/_0739_ ;
wire \myexu/myalu/_0740_ ;
wire \myexu/myalu/_0741_ ;
wire \myexu/myalu/_0742_ ;
wire \myexu/myalu/_0743_ ;
wire \myexu/myalu/_0744_ ;
wire \myexu/myalu/_0745_ ;
wire \myexu/myalu/_0746_ ;
wire \myexu/myalu/_0747_ ;
wire \myexu/myalu/_0748_ ;
wire \myexu/myalu/_0749_ ;
wire \myexu/myalu/_0750_ ;
wire \myexu/myalu/_0751_ ;
wire \myexu/myalu/_0752_ ;
wire \myexu/myalu/_0753_ ;
wire \myexu/myalu/_0754_ ;
wire \myexu/myalu/_0755_ ;
wire \myexu/myalu/_0756_ ;
wire \myexu/myalu/_0757_ ;
wire \myexu/myalu/_0758_ ;
wire \myexu/myalu/_0759_ ;
wire \myexu/myalu/_0760_ ;
wire \myexu/myalu/_0761_ ;
wire \myexu/myalu/_0762_ ;
wire \myexu/myalu/_0763_ ;
wire \myexu/myalu/_0764_ ;
wire \myexu/myalu/_0765_ ;
wire \myexu/myalu/_0766_ ;
wire \myexu/myalu/_0767_ ;
wire \myexu/myalu/_0768_ ;
wire \myexu/myalu/_0769_ ;
wire \myexu/myalu/_0770_ ;
wire \myexu/myalu/_0771_ ;
wire \myexu/myalu/_0772_ ;
wire \myexu/myalu/_0773_ ;
wire \myexu/myalu/_0774_ ;
wire \myexu/myalu/_0775_ ;
wire \myexu/myalu/_0776_ ;
wire \myexu/myalu/_0777_ ;
wire \myexu/myalu/_0778_ ;
wire \myexu/myalu/_0779_ ;
wire \myexu/myalu/_0780_ ;
wire \myexu/myalu/_0781_ ;
wire \myexu/myalu/_0782_ ;
wire \myexu/myalu/_0783_ ;
wire \myexu/myalu/_0784_ ;
wire \myexu/myalu/_0785_ ;
wire \myexu/myalu/_0786_ ;
wire \myexu/myalu/_0787_ ;
wire \myexu/myalu/_0788_ ;
wire \myexu/myalu/_0789_ ;
wire \myexu/myalu/_0790_ ;
wire \myexu/myalu/_0791_ ;
wire \myexu/myalu/_0792_ ;
wire \myexu/myalu/_0793_ ;
wire \myexu/myalu/_0794_ ;
wire \myexu/myalu/_0795_ ;
wire \myexu/myalu/_0796_ ;
wire \myexu/myalu/_0797_ ;
wire \myexu/myalu/_0798_ ;
wire \myexu/myalu/_0799_ ;
wire \myexu/myalu/_0800_ ;
wire \myexu/myalu/_0801_ ;
wire \myexu/myalu/_0802_ ;
wire \myexu/myalu/_0803_ ;
wire \myexu/myalu/_0804_ ;
wire \myexu/myalu/_0805_ ;
wire \myexu/myalu/_0806_ ;
wire \myexu/myalu/_0807_ ;
wire \myexu/myalu/_0808_ ;
wire \myexu/myalu/_0809_ ;
wire \myexu/myalu/_0810_ ;
wire \myexu/myalu/_0811_ ;
wire \myexu/myalu/_0812_ ;
wire \myexu/myalu/_0813_ ;
wire \myexu/myalu/_0814_ ;
wire \myexu/myalu/_0815_ ;
wire \myexu/myalu/_0816_ ;
wire \myexu/myalu/_0817_ ;
wire \myexu/myalu/_0818_ ;
wire \myexu/myalu/_0819_ ;
wire \myexu/myalu/_0820_ ;
wire \myexu/myalu/_0821_ ;
wire \myexu/myalu/_0822_ ;
wire \myexu/myalu/_0823_ ;
wire \myexu/myalu/_0824_ ;
wire \myexu/myalu/_0825_ ;
wire \myexu/myalu/_0826_ ;
wire \myexu/myalu/_0827_ ;
wire \myexu/myalu/_0828_ ;
wire \myexu/myalu/_0829_ ;
wire \myexu/myalu/_0830_ ;
wire \myexu/myalu/_0831_ ;
wire \myexu/myalu/_0832_ ;
wire \myexu/myalu/_0833_ ;
wire \myexu/myalu/_0834_ ;
wire \myexu/myalu/_0835_ ;
wire \myexu/myalu/_0836_ ;
wire \myexu/myalu/_0837_ ;
wire \myexu/myalu/_0838_ ;
wire \myexu/myalu/_0839_ ;
wire \myexu/myalu/_0840_ ;
wire \myexu/myalu/_0841_ ;
wire \myexu/myalu/_0842_ ;
wire \myexu/myalu/_0843_ ;
wire \myexu/myalu/_0844_ ;
wire \myexu/myalu/_0845_ ;
wire \myexu/myalu/_0846_ ;
wire \myexu/myalu/_0847_ ;
wire \myexu/myalu/_0848_ ;
wire \myexu/myalu/_0849_ ;
wire \myexu/myalu/_0850_ ;
wire \myexu/myalu/_0851_ ;
wire \myexu/myalu/_0852_ ;
wire \myexu/myalu/_0853_ ;
wire \myexu/myalu/_0854_ ;
wire \myexu/myalu/_0855_ ;
wire \myexu/myalu/_0856_ ;
wire \myexu/myalu/_0857_ ;
wire \myexu/myalu/_0858_ ;
wire \myexu/myalu/_0859_ ;
wire \myexu/myalu/_0860_ ;
wire \myexu/myalu/_0861_ ;
wire \myexu/myalu/_0862_ ;
wire \myexu/myalu/_0863_ ;
wire \myexu/myalu/_0864_ ;
wire \myexu/myalu/_0865_ ;
wire \myexu/myalu/_0866_ ;
wire \myexu/myalu/_0867_ ;
wire \myexu/myalu/_0868_ ;
wire \myexu/myalu/_0869_ ;
wire \myexu/myalu/_0870_ ;
wire \myexu/myalu/_0871_ ;
wire \myexu/myalu/_0872_ ;
wire \myexu/myalu/_0873_ ;
wire \myexu/myalu/_0874_ ;
wire \myexu/myalu/_0875_ ;
wire \myexu/myalu/_0876_ ;
wire \myexu/myalu/_0877_ ;
wire \myexu/myalu/_0878_ ;
wire \myexu/myalu/_0879_ ;
wire \myexu/myalu/_0880_ ;
wire \myexu/myalu/_0881_ ;
wire \myexu/myalu/_0882_ ;
wire \myexu/myalu/_0883_ ;
wire \myexu/myalu/_0884_ ;
wire \myexu/myalu/_0885_ ;
wire \myexu/myalu/_0886_ ;
wire \myexu/myalu/_0887_ ;
wire \myexu/myalu/_0888_ ;
wire \myexu/myalu/_0889_ ;
wire \myexu/myalu/_0890_ ;
wire \myexu/myalu/_0891_ ;
wire \myexu/myalu/_0892_ ;
wire \myexu/myalu/_0893_ ;
wire \myexu/myalu/_0894_ ;
wire \myexu/myalu/_0895_ ;
wire \myexu/myalu/_0896_ ;
wire \myexu/myalu/_0897_ ;
wire \myexu/myalu/_0898_ ;
wire \myexu/myalu/_0899_ ;
wire \myexu/myalu/_0900_ ;
wire \myexu/myalu/_0901_ ;
wire \myexu/myalu/_0902_ ;
wire \myexu/myalu/_0903_ ;
wire \myexu/myalu/_0904_ ;
wire \myexu/myalu/_0905_ ;
wire \myexu/myalu/_0906_ ;
wire \myexu/myalu/_0907_ ;
wire \myexu/myalu/_0908_ ;
wire \myexu/myalu/_0909_ ;
wire \myexu/myalu/_0910_ ;
wire \myexu/myalu/_0911_ ;
wire \myexu/myalu/_0912_ ;
wire \myexu/myalu/_0913_ ;
wire \myexu/myalu/_0914_ ;
wire \myexu/myalu/_0915_ ;
wire \myexu/myalu/_0916_ ;
wire \myexu/myalu/_0917_ ;
wire \myexu/myalu/_0918_ ;
wire \myexu/myalu/_0919_ ;
wire \myexu/myalu/_0920_ ;
wire \myexu/myalu/_0921_ ;
wire \myexu/myalu/_0922_ ;
wire \myexu/myalu/_0923_ ;
wire \myexu/myalu/_0924_ ;
wire \myexu/myalu/_0925_ ;
wire \myexu/myalu/_0926_ ;
wire \myexu/myalu/_0927_ ;
wire \myexu/myalu/_0928_ ;
wire \myexu/myalu/_0929_ ;
wire \myexu/myalu/_0930_ ;
wire \myexu/myalu/_0931_ ;
wire \myexu/myalu/_0932_ ;
wire \myexu/myalu/_0933_ ;
wire \myexu/myalu/_0934_ ;
wire \myexu/myalu/_0935_ ;
wire \myexu/myalu/_0936_ ;
wire \myexu/myalu/_0937_ ;
wire \myexu/myalu/_0938_ ;
wire \myexu/myalu/_0939_ ;
wire \myexu/myalu/_0940_ ;
wire \myexu/myalu/_0941_ ;
wire \myexu/myalu/_0942_ ;
wire \myexu/myalu/_0943_ ;
wire \myexu/myalu/_0944_ ;
wire \myexu/myalu/_0945_ ;
wire \myexu/myalu/_0946_ ;
wire \myexu/myalu/_0947_ ;
wire \myexu/myalu/_0948_ ;
wire \myexu/myalu/_0949_ ;
wire \myexu/myalu/_0950_ ;
wire \myexu/myalu/_0951_ ;
wire \myexu/myalu/_0952_ ;
wire \myexu/myalu/_0953_ ;
wire \myexu/myalu/_0954_ ;
wire \myexu/myalu/_0955_ ;
wire \myexu/myalu/_0956_ ;
wire \myexu/myalu/_0957_ ;
wire \myexu/myalu/_0958_ ;
wire \myexu/myalu/_0959_ ;
wire \myexu/myalu/_0960_ ;
wire \myexu/myalu/_0961_ ;
wire \myexu/myalu/_0962_ ;
wire \myexu/myalu/_0963_ ;
wire \myexu/myalu/_0964_ ;
wire \myexu/myalu/_0965_ ;
wire \myexu/myalu/_0966_ ;
wire \myexu/myalu/_0967_ ;
wire \myexu/myalu/_0968_ ;
wire \myexu/myalu/_0969_ ;
wire \myexu/myalu/_0970_ ;
wire \myexu/myalu/_0971_ ;
wire \myexu/myalu/_0972_ ;
wire \myexu/myalu/_0973_ ;
wire \myexu/myalu/_0974_ ;
wire \myexu/myalu/_0975_ ;
wire \myexu/myalu/_0976_ ;
wire \myexu/myalu/_0977_ ;
wire \myexu/myalu/_0978_ ;
wire \myexu/myalu/_0979_ ;
wire \myexu/myalu/_0980_ ;
wire \myexu/myalu/_0981_ ;
wire \myexu/myalu/_0982_ ;
wire \myexu/myalu/_0983_ ;
wire \myexu/myalu/_0984_ ;
wire \myexu/myalu/_0985_ ;
wire \myexu/myalu/_0986_ ;
wire \myexu/myalu/_0987_ ;
wire \myexu/myalu/_0988_ ;
wire \myexu/myalu/_0989_ ;
wire \myexu/myalu/_0990_ ;
wire \myexu/myalu/_0991_ ;
wire \myexu/myalu/_0992_ ;
wire \myexu/myalu/_0993_ ;
wire \myexu/myalu/_0994_ ;
wire \myexu/myalu/_0995_ ;
wire \myexu/myalu/_0996_ ;
wire \myexu/myalu/_0997_ ;
wire \myexu/myalu/_0998_ ;
wire \myexu/myalu/_0999_ ;
wire \myexu/myalu/_1000_ ;
wire \myexu/myalu/_1001_ ;
wire \myexu/myalu/_1002_ ;
wire \myexu/myalu/_1003_ ;
wire \myexu/myalu/_1004_ ;
wire \myexu/myalu/_1005_ ;
wire \myexu/myalu/_1006_ ;
wire \myexu/myalu/_1007_ ;
wire \myexu/myalu/_1008_ ;
wire \myexu/myalu/_1009_ ;
wire \myexu/myalu/_1010_ ;
wire \myexu/myalu/_1011_ ;
wire \myexu/myalu/_1012_ ;
wire \myexu/myalu/_1013_ ;
wire \myexu/myalu/_1014_ ;
wire \myexu/myalu/_1015_ ;
wire \myexu/myalu/_1016_ ;
wire \myexu/myalu/_1017_ ;
wire \myexu/myalu/_1018_ ;
wire \myexu/myalu/_1019_ ;
wire \myexu/myalu/_1020_ ;
wire \myexu/myalu/_1021_ ;
wire \myexu/myalu/_1022_ ;
wire \myexu/myalu/_1023_ ;
wire \myexu/myalu/_1024_ ;
wire \myexu/myalu/_1025_ ;
wire \myexu/myalu/_1026_ ;
wire \myexu/myalu/_1027_ ;
wire \myexu/myalu/_1028_ ;
wire \myexu/myalu/_1029_ ;
wire \myexu/myalu/_1030_ ;
wire \myexu/myalu/_1031_ ;
wire \myexu/myalu/_1032_ ;
wire \myexu/myalu/_1033_ ;
wire \myexu/myalu/_1034_ ;
wire \myexu/myalu/_1035_ ;
wire \myexu/myalu/_1036_ ;
wire \myexu/myalu/_1037_ ;
wire \myexu/myalu/_1038_ ;
wire \myexu/myalu/_1039_ ;
wire \myexu/myalu/_1040_ ;
wire \myexu/myalu/_1041_ ;
wire \myexu/myalu/_1042_ ;
wire \myexu/myalu/_1043_ ;
wire \myexu/myalu/_1044_ ;
wire \myexu/myalu/_1045_ ;
wire \myexu/myalu/_1046_ ;
wire \myexu/myalu/_1047_ ;
wire \myexu/myalu/_1048_ ;
wire \myexu/myalu/_1049_ ;
wire \myexu/myalu/_1050_ ;
wire \myexu/myalu/_1051_ ;
wire \myexu/myalu/_1052_ ;
wire \myexu/myalu/_1053_ ;
wire \myexu/myalu/_1054_ ;
wire \myexu/myalu/_1055_ ;
wire \myexu/myalu/_1056_ ;
wire \myexu/myalu/_1057_ ;
wire \myexu/myalu/_1058_ ;
wire \myexu/myalu/_1059_ ;
wire \myexu/myalu/_1060_ ;
wire \myexu/myalu/_1061_ ;
wire \myexu/myalu/_1062_ ;
wire \myexu/myalu/_1063_ ;
wire \myexu/myalu/_1064_ ;
wire \myexu/myalu/_1065_ ;
wire \myexu/myalu/_1066_ ;
wire \myexu/myalu/_1067_ ;
wire \myexu/myalu/_1068_ ;
wire \myexu/myalu/_1069_ ;
wire \myexu/myalu/_1070_ ;
wire \myexu/myalu/_1071_ ;
wire \myexu/myalu/_1072_ ;
wire \myexu/myalu/_1073_ ;
wire \myexu/myalu/_1074_ ;
wire \myexu/myalu/_1075_ ;
wire \myexu/myalu/_1076_ ;
wire \myexu/myalu/_1077_ ;
wire \myexu/myalu/_1078_ ;
wire \myexu/myalu/_1079_ ;
wire \myexu/myalu/_1080_ ;
wire \myexu/myalu/_1081_ ;
wire \myexu/myalu/_1082_ ;
wire \myexu/myalu/_1083_ ;
wire \myexu/myalu/_1084_ ;
wire \myexu/myalu/_1085_ ;
wire \myexu/myalu/_1086_ ;
wire \myexu/myalu/_1087_ ;
wire \myexu/myalu/_1088_ ;
wire \myexu/myalu/_1089_ ;
wire \myexu/myalu/_1090_ ;
wire \myexu/myalu/_1091_ ;
wire \myexu/myalu/_1092_ ;
wire \myexu/myalu/_1093_ ;
wire \myexu/myalu/_1094_ ;
wire \myexu/myalu/_1095_ ;
wire \myexu/myalu/_1096_ ;
wire \myexu/myalu/_1097_ ;
wire \myexu/myalu/_1098_ ;
wire \myexu/myalu/_1099_ ;
wire \myexu/myalu/_1100_ ;
wire \myexu/myalu/_1101_ ;
wire \myexu/myalu/_1102_ ;
wire \myexu/myalu/_1103_ ;
wire \myexu/myalu/_1104_ ;
wire \myexu/myalu/_1105_ ;
wire \myexu/myalu/_1106_ ;
wire \myexu/myalu/_1107_ ;
wire \myexu/myalu/_1108_ ;
wire \myexu/myalu/_1109_ ;
wire \myexu/myalu/_1110_ ;
wire \myexu/myalu/_1111_ ;
wire \myexu/myalu/_1112_ ;
wire \myexu/myalu/_1113_ ;
wire \myexu/myalu/_1114_ ;
wire \myexu/myalu/_1115_ ;
wire \myexu/myalu/_1116_ ;
wire \myexu/myalu/_1117_ ;
wire \myexu/myalu/_1118_ ;
wire \myexu/myalu/_1119_ ;
wire \myexu/myalu/_1120_ ;
wire \myexu/myalu/_1121_ ;
wire \myexu/myalu/_1122_ ;
wire \myexu/myalu/_1123_ ;
wire \myexu/myalu/_1124_ ;
wire \myexu/myalu/_1125_ ;
wire \myexu/myalu/_1126_ ;
wire \myexu/myalu/_1127_ ;
wire \myexu/myalu/_1128_ ;
wire \myexu/myalu/_1129_ ;
wire \myexu/myalu/_1130_ ;
wire \myexu/myalu/_1131_ ;
wire \myexu/myalu/_1132_ ;
wire \myexu/myalu/_1133_ ;
wire \myexu/myalu/_1134_ ;
wire \myexu/myalu/_1135_ ;
wire \myexu/myalu/_1136_ ;
wire \myexu/myalu/_1137_ ;
wire \myexu/myalu/_1138_ ;
wire \myexu/myalu/_1139_ ;
wire \myexu/myalu/_1140_ ;
wire \myexu/myalu/_1141_ ;
wire \myexu/myalu/_1142_ ;
wire \myexu/myalu/_1143_ ;
wire \myexu/myalu/_1144_ ;
wire \myexu/myalu/_1145_ ;
wire \myexu/myalu/_1146_ ;
wire \myexu/myalu/_1147_ ;
wire \myexu/myalu/_1148_ ;
wire \myexu/myalu/_1149_ ;
wire \myexu/myalu/_1150_ ;
wire \myexu/myalu/_1151_ ;
wire \myexu/myalu/_1152_ ;
wire \myexu/myalu/_1153_ ;
wire \myexu/myalu/_1154_ ;
wire \myexu/myalu/_1155_ ;
wire \myexu/myalu/_1156_ ;
wire \myexu/myalu/_1157_ ;
wire \myexu/myalu/_1158_ ;
wire \myexu/myalu/_1159_ ;
wire \myexu/myalu/_1160_ ;
wire \myexu/myalu/_1161_ ;
wire \myexu/myalu/_1162_ ;
wire \myexu/myalu/_1163_ ;
wire \myexu/myalu/_1164_ ;
wire \myexu/myalu/_1165_ ;
wire \myexu/myalu/_1166_ ;
wire \myexu/myalu/_1167_ ;
wire \myexu/myalu/_1168_ ;
wire \myexu/myalu/_1169_ ;
wire \myexu/myalu/_1170_ ;
wire \myexu/myalu/_1171_ ;
wire \myexu/myalu/_1172_ ;
wire \myexu/myalu/_1173_ ;
wire \myexu/myalu/_1174_ ;
wire \myexu/myalu/_1175_ ;
wire \myexu/myalu/_1176_ ;
wire \myexu/myalu/_1177_ ;
wire \myexu/myalu/_1178_ ;
wire \myexu/myalu/_1179_ ;
wire \myexu/myalu/_1180_ ;
wire \myexu/myalu/_1181_ ;
wire \myexu/myalu/_1182_ ;
wire \myexu/myalu/_1183_ ;
wire \myexu/myalu/_1184_ ;
wire \myexu/myalu/_1185_ ;
wire \myexu/myalu/_1186_ ;
wire \myexu/myalu/_1187_ ;
wire \myexu/myalu/_1188_ ;
wire \myexu/myalu/_1189_ ;
wire \myexu/myalu/_1190_ ;
wire \myexu/myalu/_1191_ ;
wire \myexu/myalu/_1192_ ;
wire \myexu/myalu/_1193_ ;
wire \myexu/myalu/_1194_ ;
wire \myexu/myalu/_1195_ ;
wire \myexu/myalu/_1196_ ;
wire \myexu/myalu/_1197_ ;
wire \myexu/myalu/_1198_ ;
wire \myexu/myalu/_1199_ ;
wire \myexu/myalu/_1200_ ;
wire \myexu/myalu/_1201_ ;
wire \myexu/myalu/_1202_ ;
wire \myexu/myalu/_1203_ ;
wire \myexu/myalu/_1204_ ;
wire \myexu/myalu/_1205_ ;
wire \myexu/myalu/_1206_ ;
wire \myexu/myalu/_1207_ ;
wire \myexu/myalu/_1208_ ;
wire \myexu/myalu/_1209_ ;
wire \myexu/myalu/_1210_ ;
wire \myexu/myalu/_1211_ ;
wire \myexu/myalu/_1212_ ;
wire \myexu/myalu/_1213_ ;
wire \myexu/myalu/_1214_ ;
wire \myexu/myalu/_1215_ ;
wire \myexu/myalu/_1216_ ;
wire \myexu/myalu/_1217_ ;
wire \myexu/myalu/_1218_ ;
wire \myexu/myalu/_1219_ ;
wire \myexu/myalu/_1220_ ;
wire \myexu/myalu/_1221_ ;
wire \myexu/myalu/_1222_ ;
wire \myexu/myalu/_1223_ ;
wire \myexu/myalu/_1224_ ;
wire \myexu/myalu/_1225_ ;
wire \myexu/myalu/_1226_ ;
wire \myexu/myalu/_1227_ ;
wire \myexu/myalu/_1228_ ;
wire \myexu/myalu/_1229_ ;
wire \myexu/myalu/_1230_ ;
wire \myexu/myalu/_1231_ ;
wire \myexu/myalu/_1232_ ;
wire \myexu/myalu/_1233_ ;
wire \myexu/myalu/_1234_ ;
wire \myexu/myalu/_1235_ ;
wire \myexu/myalu/_1236_ ;
wire \myexu/myalu/_1237_ ;
wire \myexu/myalu/_1238_ ;
wire \myexu/myalu/_1239_ ;
wire \myexu/myalu/_1240_ ;
wire \myexu/myalu/_1241_ ;
wire \myexu/myalu/_1242_ ;
wire \myexu/myalu/_1243_ ;
wire \myexu/myalu/_1244_ ;
wire \myexu/myalu/_1245_ ;
wire \myexu/myalu/_1246_ ;
wire \myexu/myalu/_1247_ ;
wire \myexu/myalu/_1248_ ;
wire \myexu/myalu/_1249_ ;
wire \myexu/myalu/_1250_ ;
wire \myexu/myalu/_1251_ ;
wire \myexu/myalu/_1252_ ;
wire \myexu/myalu/_1253_ ;
wire \myexu/myalu/_1254_ ;
wire \myexu/myalu/_1255_ ;
wire \myexu/myalu/_1256_ ;
wire \myexu/myalu/_1257_ ;
wire \myexu/myalu/_1258_ ;
wire \myexu/myalu/_1259_ ;
wire \myexu/myalu/_1260_ ;
wire \myexu/myalu/_1261_ ;
wire \myexu/myalu/_1262_ ;
wire \myexu/myalu/_1263_ ;
wire \myexu/myalu/_1264_ ;
wire \myexu/myalu/_1265_ ;
wire \myexu/myalu/_1266_ ;
wire \myexu/myalu/_1267_ ;
wire \myexu/myalu/_1268_ ;
wire \myexu/myalu/_1269_ ;
wire \myexu/myalu/_1270_ ;
wire \myexu/myalu/_1271_ ;
wire \myexu/myalu/_1272_ ;
wire \myexu/myalu/_1273_ ;
wire \myexu/myalu/_1274_ ;
wire \myexu/myalu/_1275_ ;
wire \myexu/myalu/_1276_ ;
wire \myexu/myalu/_1277_ ;
wire \myexu/myalu/_1278_ ;
wire \myexu/myalu/_1279_ ;
wire \myexu/myalu/_1280_ ;
wire \myexu/myalu/_1281_ ;
wire \myexu/myalu/_1282_ ;
wire \myexu/myalu/_1283_ ;
wire \myexu/myalu/_1284_ ;
wire \myexu/myalu/_1285_ ;
wire \myexu/myalu/_1286_ ;
wire \myexu/myalu/_1287_ ;
wire \myexu/myalu/_1288_ ;
wire \myexu/myalu/_1289_ ;
wire \myexu/myalu/_1290_ ;
wire \myexu/myalu/_1291_ ;
wire \myexu/myalu/_1292_ ;
wire \myexu/myalu/_1293_ ;
wire \myexu/myalu/_1294_ ;
wire \myexu/myalu/_1295_ ;
wire \myexu/myalu/_1296_ ;
wire \myexu/myalu/_1297_ ;
wire \myexu/myalu/_1298_ ;
wire \myexu/myalu/_1299_ ;
wire \myexu/myalu/_1300_ ;
wire \myexu/myalu/_1301_ ;
wire \myexu/myalu/_1302_ ;
wire \myexu/myalu/_1303_ ;
wire \myexu/myalu/_1304_ ;
wire \myexu/myalu/_1305_ ;
wire \myexu/myalu/_1306_ ;
wire \myexu/myalu/_1307_ ;
wire \myexu/myalu/_1308_ ;
wire \myexu/myalu/_1309_ ;
wire \myexu/myalu/_1310_ ;
wire \myexu/myalu/_1311_ ;
wire \myexu/myalu/_1312_ ;
wire \myexu/myalu/_1313_ ;
wire \myexu/myalu/_1314_ ;
wire \myexu/myalu/_1315_ ;
wire \myexu/myalu/_1316_ ;
wire \myexu/myalu/_1317_ ;
wire \myexu/myalu/_1318_ ;
wire \myexu/myalu/_1319_ ;
wire \myexu/myalu/_1320_ ;
wire \myexu/myalu/_1321_ ;
wire \myexu/myalu/_1322_ ;
wire \myexu/myalu/_1323_ ;
wire \myexu/myalu/_1324_ ;
wire \myexu/myalu/_1325_ ;
wire \myexu/myalu/_1326_ ;
wire \myexu/myalu/_1327_ ;
wire \myexu/myalu/_1328_ ;
wire \myexu/myalu/_1329_ ;
wire \myexu/myalu/_1330_ ;
wire \myexu/myalu/_1331_ ;
wire \myexu/myalu/_1332_ ;
wire \myexu/myalu/_1333_ ;
wire \myexu/myalu/_1334_ ;
wire \myexu/myalu/_1335_ ;
wire \myexu/myalu/_1336_ ;
wire \myexu/myalu/_1337_ ;
wire \myexu/myalu/_1338_ ;
wire \myexu/myalu/_1339_ ;
wire \myexu/myalu/_1340_ ;
wire \myexu/myalu/_1341_ ;
wire \myexu/myalu/_1342_ ;
wire \myexu/myalu/_1343_ ;
wire \myexu/myalu/_1344_ ;
wire \myexu/myalu/_1345_ ;
wire \myexu/myalu/_1346_ ;
wire \myexu/myalu/_1347_ ;
wire \myexu/myalu/_1348_ ;
wire \myexu/myalu/_1349_ ;
wire \myexu/myalu/_1350_ ;
wire \myexu/myalu/_1351_ ;
wire \myexu/myalu/_1352_ ;
wire \myexu/myalu/_1353_ ;
wire \myexu/myalu/_1354_ ;
wire \myexu/myalu/_1355_ ;
wire \myexu/myalu/_1356_ ;
wire \myexu/myalu/_1357_ ;
wire \myexu/myalu/_1358_ ;
wire \myexu/myalu/_1359_ ;
wire \myexu/myalu/_1360_ ;
wire \myexu/myalu/_1361_ ;
wire \myexu/myalu/_1362_ ;
wire \myexu/myalu/_1363_ ;
wire \myexu/myalu/_1364_ ;
wire \myexu/myalu/_1365_ ;
wire \myexu/myalu/_1366_ ;
wire \myexu/myalu/_1367_ ;
wire \myexu/myalu/_1368_ ;
wire \myexu/myalu/_1369_ ;
wire \myexu/myalu/_1370_ ;
wire \myexu/myalu/_1371_ ;
wire \myexu/myalu/_1372_ ;
wire \myexu/myalu/_1373_ ;
wire \myexu/myalu/_1374_ ;
wire \myexu/myalu/_1375_ ;
wire \myexu/myalu/_1376_ ;
wire \myexu/myalu/_1377_ ;
wire \myexu/myalu/_1378_ ;
wire \myexu/myalu/_1379_ ;
wire \myexu/myalu/_1380_ ;
wire \myexu/myalu/_1381_ ;
wire \myexu/myalu/_1382_ ;
wire \myexu/myalu/_1383_ ;
wire \myexu/myalu/_1384_ ;
wire \myexu/myalu/_1385_ ;
wire \myexu/myalu/_1386_ ;
wire \myexu/myalu/_1387_ ;
wire \myexu/myalu/_1388_ ;
wire \myexu/myalu/_1389_ ;
wire \myexu/myalu/_1390_ ;
wire \myexu/myalu/_1391_ ;
wire \myfc/_000_ ;
wire \myfc/_001_ ;
wire \myfc/_002_ ;
wire \myfc/_003_ ;
wire \myfc/_004_ ;
wire \myfc/_005_ ;
wire \myfc/_006_ ;
wire \myfc/_007_ ;
wire \myfc/_008_ ;
wire \myfc/_009_ ;
wire \myfc/_010_ ;
wire \myfc/_011_ ;
wire \myfc/_012_ ;
wire \myfc/_013_ ;
wire \myfc/_014_ ;
wire \myfc/_015_ ;
wire \myfc/_016_ ;
wire \myfc/_017_ ;
wire \myfc/_018_ ;
wire \myfc/_019_ ;
wire \myfc/_020_ ;
wire \myfc/_021_ ;
wire \myfc/_022_ ;
wire \myfc/_023_ ;
wire \myfc/_024_ ;
wire \myfc/_025_ ;
wire \myfc/_026_ ;
wire \myfc/_027_ ;
wire \myfc/_028_ ;
wire \myfc/_029_ ;
wire \myfc/_030_ ;
wire \myfc/_031_ ;
wire \myfc/_032_ ;
wire \myfc/_033_ ;
wire \myfc/_034_ ;
wire \myfc/_035_ ;
wire \myfc/_036_ ;
wire \myfc/_037_ ;
wire \myfc/_038_ ;
wire \myfc/_039_ ;
wire \myfc/_040_ ;
wire \myfc/_041_ ;
wire \myfc/_042_ ;
wire \myfc/_043_ ;
wire \myfc/_044_ ;
wire \myfc/_045_ ;
wire \myfc/_046_ ;
wire \myfc/_047_ ;
wire \myfc/_048_ ;
wire \myfc/_049_ ;
wire \myfc/_050_ ;
wire \myfc/_051_ ;
wire \myfc/_052_ ;
wire \myfc/_053_ ;
wire \myfc/_054_ ;
wire \myfc/_055_ ;
wire \myfc/_056_ ;
wire \myfc/_057_ ;
wire \myfc/_058_ ;
wire \myfc/_059_ ;
wire \myfc/_060_ ;
wire \myfc/_061_ ;
wire \myfc/_062_ ;
wire \myfc/_063_ ;
wire \myfc/_064_ ;
wire \myfc/_065_ ;
wire \myfc/_066_ ;
wire \myfc/_067_ ;
wire \myfc/_068_ ;
wire \myfc/_069_ ;
wire \myfc/_070_ ;
wire \myfc/_071_ ;
wire \myfc/_072_ ;
wire \myfc/_073_ ;
wire \myfc/_074_ ;
wire \myfc/_075_ ;
wire \myfc/_076_ ;
wire \myfc/_077_ ;
wire \myfc/_078_ ;
wire \myfc/_079_ ;
wire \myfc/_080_ ;
wire \myfc/_081_ ;
wire \myfc/_082_ ;
wire \myfc/_083_ ;
wire \myfc/_084_ ;
wire \myfc/_085_ ;
wire \myfc/_086_ ;
wire \myfc/_087_ ;
wire \myfc/_088_ ;
wire \myfc/_089_ ;
wire \myfc/_090_ ;
wire \myfc/_091_ ;
wire \myfc/_092_ ;
wire \myfc/_093_ ;
wire \myfc/_094_ ;
wire \myfc/_095_ ;
wire \myfc/_096_ ;
wire \myfc/_097_ ;
wire \myfc/_098_ ;
wire \myfc/_099_ ;
wire \myfc/_100_ ;
wire \myfc/_101_ ;
wire \myfc/_102_ ;
wire \myfc/_103_ ;
wire \myfc/_104_ ;
wire \myfc/_105_ ;
wire \myfc/_106_ ;
wire \myfc/_107_ ;
wire \myfc/_108_ ;
wire \myfc/_109_ ;
wire \myfc/_110_ ;
wire \myfc/_111_ ;
wire \myfc/_112_ ;
wire \myfc/_113_ ;
wire \myfc/_114_ ;
wire \myfc/_115_ ;
wire \myfc/_116_ ;
wire \myfc/_117_ ;
wire \myfc/_118_ ;
wire \myfc/_119_ ;
wire \myfc/_120_ ;
wire \myfc/_121_ ;
wire \myfc/_122_ ;
wire \myfc/_123_ ;
wire \myfc/_124_ ;
wire \myfc/_125_ ;
wire \myfc/_126_ ;
wire \myfc/_127_ ;
wire \myfc/_128_ ;
wire \myfc/_129_ ;
wire \myfc/_130_ ;
wire \myfc/_131_ ;
wire \myfc/_132_ ;
wire \myfc/_133_ ;
wire \myfc/_134_ ;
wire \myfc/_135_ ;
wire \myfc/_136_ ;
wire \myfc/_137_ ;
wire \myfc/_138_ ;
wire \myfc/_139_ ;
wire \myfc/_140_ ;
wire \myfc/_141_ ;
wire \myfc/_142_ ;
wire \myfc/_143_ ;
wire \myfc/_144_ ;
wire \myfc/_145_ ;
wire \myfc/_146_ ;
wire \myfc/_147_ ;
wire \myfc/_148_ ;
wire \myfc/_149_ ;
wire \myfc/_150_ ;
wire \myfc/_151_ ;
wire \myfc/_152_ ;
wire \myfc/_153_ ;
wire \myfc/_154_ ;
wire \myfc/_155_ ;
wire \myfc/_156_ ;
wire \myfc/_157_ ;
wire \myfc/_158_ ;
wire \myfc/_159_ ;
wire \myfc/_160_ ;
wire \myfc/_161_ ;
wire \myfc/_162_ ;
wire \myfc/_163_ ;
wire \myfc/_164_ ;
wire \myfc/_165_ ;
wire \myfc/_166_ ;
wire \myfc/_167_ ;
wire \myfc/_168_ ;
wire \myfc/_169_ ;
wire \myfc/_170_ ;
wire \myfc/_171_ ;
wire \myfc/_172_ ;
wire \myfc/_173_ ;
wire \myfc/_174_ ;
wire \myfc/_175_ ;
wire \myfc/_176_ ;
wire \myfc/_177_ ;
wire \myfc/_178_ ;
wire \myfc/_179_ ;
wire \myfc/_180_ ;
wire \myfc/_181_ ;
wire \myfc/_182_ ;
wire \myfc/_183_ ;
wire \myfc/_184_ ;
wire \myfc/_185_ ;
wire \myfc/_186_ ;
wire \myfc/_187_ ;
wire \myfc/_188_ ;
wire \myfc/_189_ ;
wire \myfc/_190_ ;
wire \myfc/_191_ ;
wire \myfc/_192_ ;
wire \myfc/_193_ ;
wire \myfc/_194_ ;
wire \myfc/_195_ ;
wire \myfc/_196_ ;
wire \myfc/_197_ ;
wire \myfc/_198_ ;
wire \myfc/_199_ ;
wire \myfc/_200_ ;
wire \myfc/_201_ ;
wire \myfc/_202_ ;
wire \myfc/_203_ ;
wire \myfc/_204_ ;
wire \myfc/_205_ ;
wire \myfc/_206_ ;
wire \myfc/_207_ ;
wire \myfc/_208_ ;
wire \myfc/_209_ ;
wire \myfc/_210_ ;
wire \myfc/_211_ ;
wire \myfc/_212_ ;
wire \myfc/_213_ ;
wire \myfc/_214_ ;
wire \myfc/_215_ ;
wire \myfc/_216_ ;
wire \myfc/_217_ ;
wire \myfc/_218_ ;
wire \myfc/_219_ ;
wire \myfc/_220_ ;
wire \myfc/_221_ ;
wire \myfc/_222_ ;
wire \myfc/_223_ ;
wire \myfc/_224_ ;
wire \myfc/_225_ ;
wire \myfc/_226_ ;
wire \myfc/_227_ ;
wire \myfc/_228_ ;
wire \myfc/_229_ ;
wire \myfc/_230_ ;
wire \myfc/_231_ ;
wire \myfc/_232_ ;
wire \myfc/_233_ ;
wire \myfc/_234_ ;
wire \myfc/_235_ ;
wire \myfc/_236_ ;
wire \myfc/_237_ ;
wire \myfc/_238_ ;
wire \myfc/_239_ ;
wire \myfc/_240_ ;
wire \myfc/_241_ ;
wire \myfc/_242_ ;
wire \myfc/_243_ ;
wire \myfc/_244_ ;
wire \myfc/_245_ ;
wire \myfc/_246_ ;
wire \myfc/_247_ ;
wire \myfc/_248_ ;
wire \myfc/_249_ ;
wire \myfc/_250_ ;
wire \myfc/_251_ ;
wire \myfc/_252_ ;
wire \myfc/_253_ ;
wire \myfc/_254_ ;
wire \myfc/_255_ ;
wire \myfc/_256_ ;
wire \myfc/_257_ ;
wire \myfc/_258_ ;
wire \myfc/_259_ ;
wire \myfc/_260_ ;
wire \myfc/_261_ ;
wire \myfc/_262_ ;
wire \myfc/_263_ ;
wire \myfc/_264_ ;
wire \myfc/_265_ ;
wire \myfc/_266_ ;
wire \myfc/_267_ ;
wire \myfc/_268_ ;
wire \myfc/_269_ ;
wire \myfc/_270_ ;
wire \myfc/_271_ ;
wire \myfc/_272_ ;
wire \myfc/_273_ ;
wire \myfc/_274_ ;
wire \myfc/_275_ ;
wire \myfc/_276_ ;
wire \myfc/_277_ ;
wire \myfc/_278_ ;
wire \myfc/_279_ ;
wire \myfc/_280_ ;
wire \myfc/_281_ ;
wire \myfc/_282_ ;
wire \myfc/_283_ ;
wire \myfc/_284_ ;
wire \myfc/_285_ ;
wire \myfc/_286_ ;
wire \myfc/_287_ ;
wire \myfc/_288_ ;
wire \myfc/_289_ ;
wire \myfc/_290_ ;
wire \myfc/_291_ ;
wire \myfc/_292_ ;
wire \myfc/_293_ ;
wire \myfc/_294_ ;
wire \myfc/_295_ ;
wire \myfc/_296_ ;
wire \myfc/_297_ ;
wire \myfc/_298_ ;
wire \myfc/_299_ ;
wire \myfc/_300_ ;
wire \myfc/_301_ ;
wire \myfc/_302_ ;
wire \myfc/_303_ ;
wire \myfc/_304_ ;
wire \myfc/_305_ ;
wire \myfc/_306_ ;
wire \myfc/_307_ ;
wire \myfc/_308_ ;
wire \myfc/_309_ ;
wire \myfc/_310_ ;
wire \myfc/_311_ ;
wire \myfc/_312_ ;
wire \myfc/_313_ ;
wire \myfc/_314_ ;
wire \myfc/_315_ ;
wire \myfc/_316_ ;
wire \myfc/_317_ ;
wire \myfc/_318_ ;
wire \myfc/_319_ ;
wire \myfc/_320_ ;
wire \myfc/_321_ ;
wire \myfc/_322_ ;
wire \myfc/_323_ ;
wire \myfc/_324_ ;
wire \myfc/_325_ ;
wire \myfc/_326_ ;
wire \myfc/_327_ ;
wire \myfc/_328_ ;
wire \myfc/_329_ ;
wire \myfc/_330_ ;
wire \myfc/_331_ ;
wire \myfc/_332_ ;
wire \myfc/_333_ ;
wire \myfc/_334_ ;
wire \myfc/_335_ ;
wire \myfc/_336_ ;
wire \myfc/_337_ ;
wire \myfc/_338_ ;
wire \myfc/_339_ ;
wire \myfc/_340_ ;
wire \myfc/_341_ ;
wire \myfc/_342_ ;
wire \myfc/_343_ ;
wire \myfc/_344_ ;
wire \myfc/_345_ ;
wire \myfc/_346_ ;
wire \myfc/_347_ ;
wire \myfc/_348_ ;
wire \myfc/_349_ ;
wire \myfc/_350_ ;
wire \myfc/_351_ ;
wire \myfc/_352_ ;
wire \myfc/_353_ ;
wire \myfc/_354_ ;
wire \myfc/_355_ ;
wire \myfc/_356_ ;
wire \myfc/_357_ ;
wire \myfc/_358_ ;
wire \myfc/_359_ ;
wire \myfc/_360_ ;
wire \myfc/_361_ ;
wire \myfc/_362_ ;
wire \myfc/_363_ ;
wire \myfc/_364_ ;
wire \myfc/_365_ ;
wire \myfc/_366_ ;
wire \myfc/_367_ ;
wire \myfc/_368_ ;
wire \myfc/_369_ ;
wire \myfc/_370_ ;
wire \myfc/_371_ ;
wire \myfc/_372_ ;
wire \myfc/_373_ ;
wire \myfc/_374_ ;
wire \myfc/_375_ ;
wire \myfc/_376_ ;
wire \myfc/_377_ ;
wire \myfc/_378_ ;
wire \myfc/_379_ ;
wire \myfc/_380_ ;
wire \myfc/_381_ ;
wire \myfc/_382_ ;
wire \myfc/_383_ ;
wire \myfc/_384_ ;
wire \myidu/_0000_ ;
wire \myidu/_0001_ ;
wire \myidu/_0002_ ;
wire \myidu/_0003_ ;
wire \myidu/_0004_ ;
wire \myidu/_0005_ ;
wire \myidu/_0006_ ;
wire \myidu/_0007_ ;
wire \myidu/_0008_ ;
wire \myidu/_0009_ ;
wire \myidu/_0010_ ;
wire \myidu/_0011_ ;
wire \myidu/_0012_ ;
wire \myidu/_0013_ ;
wire \myidu/_0014_ ;
wire \myidu/_0015_ ;
wire \myidu/_0016_ ;
wire \myidu/_0017_ ;
wire \myidu/_0018_ ;
wire \myidu/_0019_ ;
wire \myidu/_0020_ ;
wire \myidu/_0021_ ;
wire \myidu/_0022_ ;
wire \myidu/_0023_ ;
wire \myidu/_0024_ ;
wire \myidu/_0025_ ;
wire \myidu/_0026_ ;
wire \myidu/_0027_ ;
wire \myidu/_0028_ ;
wire \myidu/_0029_ ;
wire \myidu/_0030_ ;
wire \myidu/_0031_ ;
wire \myidu/_0032_ ;
wire \myidu/_0033_ ;
wire \myidu/_0034_ ;
wire \myidu/_0035_ ;
wire \myidu/_0036_ ;
wire \myidu/_0037_ ;
wire \myidu/_0038_ ;
wire \myidu/_0039_ ;
wire \myidu/_0040_ ;
wire \myidu/_0041_ ;
wire \myidu/_0042_ ;
wire \myidu/_0043_ ;
wire \myidu/_0044_ ;
wire \myidu/_0045_ ;
wire \myidu/_0046_ ;
wire \myidu/_0047_ ;
wire \myidu/_0048_ ;
wire \myidu/_0049_ ;
wire \myidu/_0050_ ;
wire \myidu/_0051_ ;
wire \myidu/_0052_ ;
wire \myidu/_0053_ ;
wire \myidu/_0054_ ;
wire \myidu/_0055_ ;
wire \myidu/_0056_ ;
wire \myidu/_0057_ ;
wire \myidu/_0058_ ;
wire \myidu/_0059_ ;
wire \myidu/_0060_ ;
wire \myidu/_0061_ ;
wire \myidu/_0062_ ;
wire \myidu/_0063_ ;
wire \myidu/_0064_ ;
wire \myidu/_0065_ ;
wire \myidu/_0066_ ;
wire \myidu/_0067_ ;
wire \myidu/_0068_ ;
wire \myidu/_0069_ ;
wire \myidu/_0070_ ;
wire \myidu/_0071_ ;
wire \myidu/_0072_ ;
wire \myidu/_0073_ ;
wire \myidu/_0074_ ;
wire \myidu/_0075_ ;
wire \myidu/_0076_ ;
wire \myidu/_0077_ ;
wire \myidu/_0078_ ;
wire \myidu/_0079_ ;
wire \myidu/_0080_ ;
wire \myidu/_0081_ ;
wire \myidu/_0082_ ;
wire \myidu/_0083_ ;
wire \myidu/_0084_ ;
wire \myidu/_0085_ ;
wire \myidu/_0086_ ;
wire \myidu/_0087_ ;
wire \myidu/_0088_ ;
wire \myidu/_0089_ ;
wire \myidu/_0090_ ;
wire \myidu/_0091_ ;
wire \myidu/_0092_ ;
wire \myidu/_0093_ ;
wire \myidu/_0094_ ;
wire \myidu/_0095_ ;
wire \myidu/_0096_ ;
wire \myidu/_0097_ ;
wire \myidu/_0098_ ;
wire \myidu/_0099_ ;
wire \myidu/_0100_ ;
wire \myidu/_0101_ ;
wire \myidu/_0102_ ;
wire \myidu/_0103_ ;
wire \myidu/_0104_ ;
wire \myidu/_0105_ ;
wire \myidu/_0106_ ;
wire \myidu/_0107_ ;
wire \myidu/_0108_ ;
wire \myidu/_0109_ ;
wire \myidu/_0110_ ;
wire \myidu/_0111_ ;
wire \myidu/_0112_ ;
wire \myidu/_0113_ ;
wire \myidu/_0114_ ;
wire \myidu/_0115_ ;
wire \myidu/_0116_ ;
wire \myidu/_0117_ ;
wire \myidu/_0118_ ;
wire \myidu/_0119_ ;
wire \myidu/_0120_ ;
wire \myidu/_0121_ ;
wire \myidu/_0122_ ;
wire \myidu/_0123_ ;
wire \myidu/_0124_ ;
wire \myidu/_0125_ ;
wire \myidu/_0126_ ;
wire \myidu/_0127_ ;
wire \myidu/_0128_ ;
wire \myidu/_0129_ ;
wire \myidu/_0130_ ;
wire \myidu/_0131_ ;
wire \myidu/_0132_ ;
wire \myidu/_0133_ ;
wire \myidu/_0134_ ;
wire \myidu/_0135_ ;
wire \myidu/_0136_ ;
wire \myidu/_0137_ ;
wire \myidu/_0138_ ;
wire \myidu/_0139_ ;
wire \myidu/_0140_ ;
wire \myidu/_0141_ ;
wire \myidu/_0142_ ;
wire \myidu/_0143_ ;
wire \myidu/_0144_ ;
wire \myidu/_0145_ ;
wire \myidu/_0146_ ;
wire \myidu/_0147_ ;
wire \myidu/_0148_ ;
wire \myidu/_0149_ ;
wire \myidu/_0150_ ;
wire \myidu/_0151_ ;
wire \myidu/_0152_ ;
wire \myidu/_0153_ ;
wire \myidu/_0154_ ;
wire \myidu/_0155_ ;
wire \myidu/_0156_ ;
wire \myidu/_0157_ ;
wire \myidu/_0158_ ;
wire \myidu/_0159_ ;
wire \myidu/_0160_ ;
wire \myidu/_0161_ ;
wire \myidu/_0162_ ;
wire \myidu/_0163_ ;
wire \myidu/_0164_ ;
wire \myidu/_0165_ ;
wire \myidu/_0166_ ;
wire \myidu/_0167_ ;
wire \myidu/_0168_ ;
wire \myidu/_0169_ ;
wire \myidu/_0170_ ;
wire \myidu/_0171_ ;
wire \myidu/_0172_ ;
wire \myidu/_0173_ ;
wire \myidu/_0174_ ;
wire \myidu/_0175_ ;
wire \myidu/_0176_ ;
wire \myidu/_0177_ ;
wire \myidu/_0178_ ;
wire \myidu/_0179_ ;
wire \myidu/_0180_ ;
wire \myidu/_0181_ ;
wire \myidu/_0182_ ;
wire \myidu/_0183_ ;
wire \myidu/_0184_ ;
wire \myidu/_0185_ ;
wire \myidu/_0186_ ;
wire \myidu/_0187_ ;
wire \myidu/_0188_ ;
wire \myidu/_0189_ ;
wire \myidu/_0190_ ;
wire \myidu/_0191_ ;
wire \myidu/_0192_ ;
wire \myidu/_0193_ ;
wire \myidu/_0194_ ;
wire \myidu/_0195_ ;
wire \myidu/_0196_ ;
wire \myidu/_0197_ ;
wire \myidu/_0198_ ;
wire \myidu/_0199_ ;
wire \myidu/_0200_ ;
wire \myidu/_0201_ ;
wire \myidu/_0202_ ;
wire \myidu/_0203_ ;
wire \myidu/_0204_ ;
wire \myidu/_0205_ ;
wire \myidu/_0206_ ;
wire \myidu/_0207_ ;
wire \myidu/_0208_ ;
wire \myidu/_0209_ ;
wire \myidu/_0210_ ;
wire \myidu/_0211_ ;
wire \myidu/_0212_ ;
wire \myidu/_0213_ ;
wire \myidu/_0214_ ;
wire \myidu/_0215_ ;
wire \myidu/_0216_ ;
wire \myidu/_0217_ ;
wire \myidu/_0218_ ;
wire \myidu/_0219_ ;
wire \myidu/_0220_ ;
wire \myidu/_0221_ ;
wire \myidu/_0222_ ;
wire \myidu/_0223_ ;
wire \myidu/_0224_ ;
wire \myidu/_0225_ ;
wire \myidu/_0226_ ;
wire \myidu/_0227_ ;
wire \myidu/_0228_ ;
wire \myidu/_0229_ ;
wire \myidu/_0230_ ;
wire \myidu/_0231_ ;
wire \myidu/_0232_ ;
wire \myidu/_0233_ ;
wire \myidu/_0234_ ;
wire \myidu/_0235_ ;
wire \myidu/_0236_ ;
wire \myidu/_0237_ ;
wire \myidu/_0238_ ;
wire \myidu/_0239_ ;
wire \myidu/_0240_ ;
wire \myidu/_0241_ ;
wire \myidu/_0242_ ;
wire \myidu/_0243_ ;
wire \myidu/_0244_ ;
wire \myidu/_0245_ ;
wire \myidu/_0246_ ;
wire \myidu/_0247_ ;
wire \myidu/_0248_ ;
wire \myidu/_0249_ ;
wire \myidu/_0250_ ;
wire \myidu/_0251_ ;
wire \myidu/_0252_ ;
wire \myidu/_0253_ ;
wire \myidu/_0254_ ;
wire \myidu/_0255_ ;
wire \myidu/_0256_ ;
wire \myidu/_0257_ ;
wire \myidu/_0258_ ;
wire \myidu/_0259_ ;
wire \myidu/_0260_ ;
wire \myidu/_0261_ ;
wire \myidu/_0262_ ;
wire \myidu/_0263_ ;
wire \myidu/_0264_ ;
wire \myidu/_0265_ ;
wire \myidu/_0266_ ;
wire \myidu/_0267_ ;
wire \myidu/_0268_ ;
wire \myidu/_0269_ ;
wire \myidu/_0270_ ;
wire \myidu/_0271_ ;
wire \myidu/_0272_ ;
wire \myidu/_0273_ ;
wire \myidu/_0274_ ;
wire \myidu/_0275_ ;
wire \myidu/_0276_ ;
wire \myidu/_0277_ ;
wire \myidu/_0278_ ;
wire \myidu/_0279_ ;
wire \myidu/_0280_ ;
wire \myidu/_0281_ ;
wire \myidu/_0282_ ;
wire \myidu/_0283_ ;
wire \myidu/_0284_ ;
wire \myidu/_0285_ ;
wire \myidu/_0286_ ;
wire \myidu/_0287_ ;
wire \myidu/_0288_ ;
wire \myidu/_0289_ ;
wire \myidu/_0290_ ;
wire \myidu/_0291_ ;
wire \myidu/_0292_ ;
wire \myidu/_0293_ ;
wire \myidu/_0294_ ;
wire \myidu/_0295_ ;
wire \myidu/_0296_ ;
wire \myidu/_0297_ ;
wire \myidu/_0298_ ;
wire \myidu/_0299_ ;
wire \myidu/_0300_ ;
wire \myidu/_0301_ ;
wire \myidu/_0302_ ;
wire \myidu/_0303_ ;
wire \myidu/_0304_ ;
wire \myidu/_0305_ ;
wire \myidu/_0306_ ;
wire \myidu/_0307_ ;
wire \myidu/_0308_ ;
wire \myidu/_0309_ ;
wire \myidu/_0310_ ;
wire \myidu/_0311_ ;
wire \myidu/_0312_ ;
wire \myidu/_0313_ ;
wire \myidu/_0314_ ;
wire \myidu/_0315_ ;
wire \myidu/_0316_ ;
wire \myidu/_0317_ ;
wire \myidu/_0318_ ;
wire \myidu/_0319_ ;
wire \myidu/_0320_ ;
wire \myidu/_0321_ ;
wire \myidu/_0322_ ;
wire \myidu/_0323_ ;
wire \myidu/_0324_ ;
wire \myidu/_0325_ ;
wire \myidu/_0326_ ;
wire \myidu/_0327_ ;
wire \myidu/_0328_ ;
wire \myidu/_0329_ ;
wire \myidu/_0330_ ;
wire \myidu/_0331_ ;
wire \myidu/_0332_ ;
wire \myidu/_0333_ ;
wire \myidu/_0334_ ;
wire \myidu/_0335_ ;
wire \myidu/_0336_ ;
wire \myidu/_0337_ ;
wire \myidu/_0338_ ;
wire \myidu/_0339_ ;
wire \myidu/_0340_ ;
wire \myidu/_0341_ ;
wire \myidu/_0342_ ;
wire \myidu/_0343_ ;
wire \myidu/_0344_ ;
wire \myidu/_0345_ ;
wire \myidu/_0346_ ;
wire \myidu/_0347_ ;
wire \myidu/_0348_ ;
wire \myidu/_0349_ ;
wire \myidu/_0350_ ;
wire \myidu/_0351_ ;
wire \myidu/_0352_ ;
wire \myidu/_0353_ ;
wire \myidu/_0354_ ;
wire \myidu/_0355_ ;
wire \myidu/_0356_ ;
wire \myidu/_0357_ ;
wire \myidu/_0358_ ;
wire \myidu/_0359_ ;
wire \myidu/_0360_ ;
wire \myidu/_0361_ ;
wire \myidu/_0362_ ;
wire \myidu/_0363_ ;
wire \myidu/_0364_ ;
wire \myidu/_0365_ ;
wire \myidu/_0366_ ;
wire \myidu/_0367_ ;
wire \myidu/_0368_ ;
wire \myidu/_0369_ ;
wire \myidu/_0370_ ;
wire \myidu/_0371_ ;
wire \myidu/_0372_ ;
wire \myidu/_0373_ ;
wire \myidu/_0374_ ;
wire \myidu/_0375_ ;
wire \myidu/_0376_ ;
wire \myidu/_0377_ ;
wire \myidu/_0378_ ;
wire \myidu/_0379_ ;
wire \myidu/_0380_ ;
wire \myidu/_0381_ ;
wire \myidu/_0382_ ;
wire \myidu/_0383_ ;
wire \myidu/_0384_ ;
wire \myidu/_0385_ ;
wire \myidu/_0386_ ;
wire \myidu/_0387_ ;
wire \myidu/_0388_ ;
wire \myidu/_0389_ ;
wire \myidu/_0390_ ;
wire \myidu/_0391_ ;
wire \myidu/_0392_ ;
wire \myidu/_0393_ ;
wire \myidu/_0394_ ;
wire \myidu/_0395_ ;
wire \myidu/_0396_ ;
wire \myidu/_0397_ ;
wire \myidu/_0398_ ;
wire \myidu/_0399_ ;
wire \myidu/_0400_ ;
wire \myidu/_0401_ ;
wire \myidu/_0402_ ;
wire \myidu/_0403_ ;
wire \myidu/_0404_ ;
wire \myidu/_0405_ ;
wire \myidu/_0406_ ;
wire \myidu/_0407_ ;
wire \myidu/_0408_ ;
wire \myidu/_0409_ ;
wire \myidu/_0410_ ;
wire \myidu/_0411_ ;
wire \myidu/_0412_ ;
wire \myidu/_0413_ ;
wire \myidu/_0414_ ;
wire \myidu/_0415_ ;
wire \myidu/_0416_ ;
wire \myidu/_0417_ ;
wire \myidu/_0418_ ;
wire \myidu/_0419_ ;
wire \myidu/_0420_ ;
wire \myidu/_0421_ ;
wire \myidu/_0422_ ;
wire \myidu/_0423_ ;
wire \myidu/_0424_ ;
wire \myidu/_0425_ ;
wire \myidu/_0426_ ;
wire \myidu/_0427_ ;
wire \myidu/_0428_ ;
wire \myidu/_0429_ ;
wire \myidu/_0430_ ;
wire \myidu/_0431_ ;
wire \myidu/_0432_ ;
wire \myidu/_0433_ ;
wire \myidu/_0434_ ;
wire \myidu/_0435_ ;
wire \myidu/_0436_ ;
wire \myidu/_0437_ ;
wire \myidu/_0438_ ;
wire \myidu/_0439_ ;
wire \myidu/_0440_ ;
wire \myidu/_0441_ ;
wire \myidu/_0442_ ;
wire \myidu/_0443_ ;
wire \myidu/_0444_ ;
wire \myidu/_0445_ ;
wire \myidu/_0446_ ;
wire \myidu/_0447_ ;
wire \myidu/_0448_ ;
wire \myidu/_0449_ ;
wire \myidu/_0450_ ;
wire \myidu/_0451_ ;
wire \myidu/_0452_ ;
wire \myidu/_0453_ ;
wire \myidu/_0454_ ;
wire \myidu/_0455_ ;
wire \myidu/_0456_ ;
wire \myidu/_0457_ ;
wire \myidu/_0458_ ;
wire \myidu/_0459_ ;
wire \myidu/_0460_ ;
wire \myidu/_0461_ ;
wire \myidu/_0462_ ;
wire \myidu/_0463_ ;
wire \myidu/_0464_ ;
wire \myidu/_0465_ ;
wire \myidu/_0466_ ;
wire \myidu/_0467_ ;
wire \myidu/_0468_ ;
wire \myidu/_0469_ ;
wire \myidu/_0470_ ;
wire \myidu/_0471_ ;
wire \myidu/_0472_ ;
wire \myidu/_0473_ ;
wire \myidu/_0474_ ;
wire \myidu/_0475_ ;
wire \myidu/_0476_ ;
wire \myidu/_0477_ ;
wire \myidu/_0478_ ;
wire \myidu/_0479_ ;
wire \myidu/_0480_ ;
wire \myidu/_0481_ ;
wire \myidu/_0482_ ;
wire \myidu/_0483_ ;
wire \myidu/_0484_ ;
wire \myidu/_0485_ ;
wire \myidu/_0486_ ;
wire \myidu/_0487_ ;
wire \myidu/_0488_ ;
wire \myidu/_0489_ ;
wire \myidu/_0490_ ;
wire \myidu/_0491_ ;
wire \myidu/_0492_ ;
wire \myidu/_0493_ ;
wire \myidu/_0494_ ;
wire \myidu/_0495_ ;
wire \myidu/_0496_ ;
wire \myidu/_0497_ ;
wire \myidu/_0498_ ;
wire \myidu/_0499_ ;
wire \myidu/_0500_ ;
wire \myidu/_0501_ ;
wire \myidu/_0502_ ;
wire \myidu/_0503_ ;
wire \myidu/_0504_ ;
wire \myidu/_0505_ ;
wire \myidu/_0506_ ;
wire \myidu/_0507_ ;
wire \myidu/_0508_ ;
wire \myidu/_0509_ ;
wire \myidu/_0510_ ;
wire \myidu/_0511_ ;
wire \myidu/_0512_ ;
wire \myidu/_0513_ ;
wire \myidu/_0514_ ;
wire \myidu/_0515_ ;
wire \myidu/_0516_ ;
wire \myidu/_0517_ ;
wire \myidu/_0518_ ;
wire \myidu/_0519_ ;
wire \myidu/_0520_ ;
wire \myidu/_0521_ ;
wire \myidu/_0522_ ;
wire \myidu/_0523_ ;
wire \myidu/_0524_ ;
wire \myidu/_0525_ ;
wire \myidu/_0526_ ;
wire \myidu/_0527_ ;
wire \myidu/_0528_ ;
wire \myidu/_0529_ ;
wire \myidu/_0530_ ;
wire \myidu/_0531_ ;
wire \myidu/_0532_ ;
wire \myidu/_0533_ ;
wire \myidu/_0534_ ;
wire \myidu/_0535_ ;
wire \myidu/_0536_ ;
wire \myidu/_0537_ ;
wire \myidu/_0538_ ;
wire \myidu/_0539_ ;
wire \myidu/_0540_ ;
wire \myidu/_0541_ ;
wire \myidu/_0542_ ;
wire \myidu/_0543_ ;
wire \myidu/_0544_ ;
wire \myidu/_0545_ ;
wire \myidu/_0546_ ;
wire \myidu/_0547_ ;
wire \myidu/_0548_ ;
wire \myidu/_0549_ ;
wire \myidu/_0550_ ;
wire \myidu/_0551_ ;
wire \myidu/_0552_ ;
wire \myidu/_0553_ ;
wire \myidu/_0554_ ;
wire \myidu/_0555_ ;
wire \myidu/_0556_ ;
wire \myidu/_0557_ ;
wire \myidu/_0558_ ;
wire \myidu/_0559_ ;
wire \myidu/_0560_ ;
wire \myidu/_0561_ ;
wire \myidu/_0562_ ;
wire \myidu/_0563_ ;
wire \myidu/_0564_ ;
wire \myidu/_0565_ ;
wire \myidu/_0566_ ;
wire \myidu/_0567_ ;
wire \myidu/_0568_ ;
wire \myidu/_0569_ ;
wire \myidu/_0570_ ;
wire \myidu/_0571_ ;
wire \myidu/_0572_ ;
wire \myidu/_0573_ ;
wire \myidu/_0574_ ;
wire \myidu/_0575_ ;
wire \myidu/_0576_ ;
wire \myidu/_0577_ ;
wire \myidu/_0578_ ;
wire \myidu/_0579_ ;
wire \myidu/_0580_ ;
wire \myidu/_0581_ ;
wire \myidu/_0582_ ;
wire \myidu/_0583_ ;
wire \myidu/_0584_ ;
wire \myidu/_0585_ ;
wire \myidu/_0586_ ;
wire \myidu/_0587_ ;
wire \myidu/_0588_ ;
wire \myidu/_0589_ ;
wire \myidu/_0590_ ;
wire \myidu/_0591_ ;
wire \myidu/_0592_ ;
wire \myidu/_0593_ ;
wire \myidu/_0594_ ;
wire \myidu/_0595_ ;
wire \myidu/_0596_ ;
wire \myidu/_0597_ ;
wire \myidu/_0598_ ;
wire \myidu/_0599_ ;
wire \myidu/_0600_ ;
wire \myidu/_0601_ ;
wire \myidu/_0602_ ;
wire \myidu/_0603_ ;
wire \myidu/_0604_ ;
wire \myidu/_0605_ ;
wire \myidu/_0606_ ;
wire \myidu/_0607_ ;
wire \myidu/_0608_ ;
wire \myidu/_0609_ ;
wire \myidu/_0610_ ;
wire \myidu/_0611_ ;
wire \myidu/_0612_ ;
wire \myidu/_0613_ ;
wire \myidu/_0614_ ;
wire \myidu/_0615_ ;
wire \myidu/_0616_ ;
wire \myidu/_0617_ ;
wire \myidu/_0618_ ;
wire \myidu/_0619_ ;
wire \myidu/_0620_ ;
wire \myidu/_0621_ ;
wire \myidu/_0622_ ;
wire \myidu/_0623_ ;
wire \myidu/_0624_ ;
wire \myidu/_0625_ ;
wire \myidu/_0626_ ;
wire \myidu/_0627_ ;
wire \myidu/_0628_ ;
wire \myidu/_0629_ ;
wire \myidu/_0630_ ;
wire \myidu/_0631_ ;
wire \myidu/_0632_ ;
wire \myidu/_0633_ ;
wire \myidu/_0634_ ;
wire \myidu/_0635_ ;
wire \myidu/_0636_ ;
wire \myidu/_0637_ ;
wire \myidu/_0638_ ;
wire \myidu/_0639_ ;
wire \myidu/_0640_ ;
wire \myidu/_0641_ ;
wire \myidu/_0642_ ;
wire \myidu/_0643_ ;
wire \myidu/_0644_ ;
wire \myidu/_0645_ ;
wire \myidu/_0646_ ;
wire \myidu/_0647_ ;
wire \myidu/_0648_ ;
wire \myidu/_0649_ ;
wire \myidu/_0650_ ;
wire \myidu/_0651_ ;
wire \myidu/_0652_ ;
wire \myidu/_0653_ ;
wire \myidu/_0654_ ;
wire \myidu/_0655_ ;
wire \myidu/_0656_ ;
wire \myidu/_0657_ ;
wire \myidu/_0658_ ;
wire \myidu/_0659_ ;
wire \myidu/_0660_ ;
wire \myidu/_0661_ ;
wire \myidu/_0662_ ;
wire \myidu/_0663_ ;
wire \myidu/_0664_ ;
wire \myidu/_0665_ ;
wire \myidu/_0666_ ;
wire \myidu/_0667_ ;
wire \myidu/_0668_ ;
wire \myidu/_0669_ ;
wire \myidu/_0670_ ;
wire \myidu/_0671_ ;
wire \myidu/_0672_ ;
wire \myidu/_0673_ ;
wire \myidu/_0674_ ;
wire \myidu/_0675_ ;
wire \myidu/_0676_ ;
wire \myidu/_0677_ ;
wire \myidu/_0678_ ;
wire \myidu/_0679_ ;
wire \myidu/_0680_ ;
wire \myidu/_0681_ ;
wire \myidu/_0682_ ;
wire \myidu/_0683_ ;
wire \myidu/_0684_ ;
wire \myidu/_0685_ ;
wire \myidu/_0686_ ;
wire \myidu/_0687_ ;
wire \myidu/_0688_ ;
wire \myidu/_0689_ ;
wire \myidu/_0690_ ;
wire \myidu/_0691_ ;
wire \myidu/_0692_ ;
wire \myidu/_0693_ ;
wire \myidu/_0694_ ;
wire \myidu/_0695_ ;
wire \myidu/_0696_ ;
wire \myidu/_0697_ ;
wire \myidu/_0698_ ;
wire \myidu/_0699_ ;
wire \myidu/_0700_ ;
wire \myidu/_0701_ ;
wire \myidu/_0702_ ;
wire \myidu/_0703_ ;
wire \myidu/_0704_ ;
wire \myidu/_0705_ ;
wire \myidu/_0706_ ;
wire \myidu/_0707_ ;
wire \myidu/_0708_ ;
wire \myidu/_0709_ ;
wire \myidu/_0710_ ;
wire \myidu/_0711_ ;
wire \myidu/_0712_ ;
wire \myidu/_0713_ ;
wire \myidu/_0714_ ;
wire \myidu/_0715_ ;
wire \myidu/_0716_ ;
wire \myidu/_0717_ ;
wire \myidu/_0718_ ;
wire \myidu/_0719_ ;
wire \myidu/_0720_ ;
wire \myidu/_0721_ ;
wire \myidu/_0722_ ;
wire \myidu/_0723_ ;
wire \myidu/_0724_ ;
wire \myidu/_0725_ ;
wire \myidu/_0726_ ;
wire \myidu/_0727_ ;
wire \myidu/_0728_ ;
wire \myidu/_0729_ ;
wire \myidu/_0730_ ;
wire \myidu/_0731_ ;
wire \myidu/_0732_ ;
wire \myidu/_0733_ ;
wire \myidu/_0734_ ;
wire \myidu/_0735_ ;
wire \myidu/_0736_ ;
wire \myidu/_0737_ ;
wire \myidu/_0738_ ;
wire \myidu/_0739_ ;
wire \myidu/_0740_ ;
wire \myidu/_0741_ ;
wire \myidu/_0742_ ;
wire \myidu/_0743_ ;
wire \myidu/_0744_ ;
wire \myidu/_0745_ ;
wire \myidu/_0746_ ;
wire \myidu/_0747_ ;
wire \myidu/_0748_ ;
wire \myidu/_0749_ ;
wire \myidu/_0750_ ;
wire \myidu/_0751_ ;
wire \myidu/_0752_ ;
wire \myidu/_0753_ ;
wire \myidu/_0754_ ;
wire \myidu/_0755_ ;
wire \myidu/_0756_ ;
wire \myidu/_0757_ ;
wire \myidu/_0758_ ;
wire \myidu/_0759_ ;
wire \myidu/_0760_ ;
wire \myidu/_0761_ ;
wire \myidu/_0762_ ;
wire \myidu/_0763_ ;
wire \myidu/_0764_ ;
wire \myidu/_0765_ ;
wire \myidu/_0766_ ;
wire \myidu/_0767_ ;
wire \myidu/_0768_ ;
wire \myidu/_0769_ ;
wire \myidu/_0770_ ;
wire \myidu/_0771_ ;
wire \myidu/_0772_ ;
wire \myidu/_0773_ ;
wire \myidu/_0774_ ;
wire \myidu/_0775_ ;
wire \myidu/_0776_ ;
wire \myidu/_0777_ ;
wire \myidu/_0778_ ;
wire \myidu/_0779_ ;
wire \myidu/_0780_ ;
wire \myidu/_0781_ ;
wire \myidu/_0782_ ;
wire \myidu/_0783_ ;
wire \myidu/_0784_ ;
wire \myidu/_0785_ ;
wire \myidu/_0786_ ;
wire \myidu/_0787_ ;
wire \myidu/_0788_ ;
wire \myidu/_0789_ ;
wire \myidu/_0790_ ;
wire \myidu/_0791_ ;
wire \myidu/_0792_ ;
wire \myidu/_0793_ ;
wire \myidu/_0794_ ;
wire \myidu/_0795_ ;
wire \myidu/_0796_ ;
wire \myidu/_0797_ ;
wire \myidu/_0798_ ;
wire \myidu/_0799_ ;
wire \myidu/_0800_ ;
wire \myidu/_0801_ ;
wire \myidu/_0802_ ;
wire \myidu/_0803_ ;
wire \myidu/_0804_ ;
wire \myidu/_0805_ ;
wire \myidu/_0806_ ;
wire \myidu/_0807_ ;
wire \myidu/_0808_ ;
wire \myidu/_0809_ ;
wire \myidu/_0810_ ;
wire \myidu/_0811_ ;
wire \myidu/_0812_ ;
wire \myidu/_0813_ ;
wire \myidu/_0814_ ;
wire \myidu/_0815_ ;
wire \myidu/_0816_ ;
wire \myidu/_0817_ ;
wire \myidu/_0818_ ;
wire \myidu/_0819_ ;
wire \myidu/_0820_ ;
wire \myidu/_0821_ ;
wire \myidu/_0822_ ;
wire \myidu/_0823_ ;
wire \myidu/_0824_ ;
wire \myidu/_0825_ ;
wire \myidu/_0826_ ;
wire \myidu/_0827_ ;
wire \myidu/_0828_ ;
wire \myidu/_0829_ ;
wire \myidu/_0830_ ;
wire \myidu/_0831_ ;
wire \myidu/_0832_ ;
wire \myidu/_0833_ ;
wire \myidu/_0834_ ;
wire \myidu/_0835_ ;
wire \myidu/_0836_ ;
wire \myidu/_0837_ ;
wire \myidu/_0838_ ;
wire \myidu/_0839_ ;
wire \myidu/_0840_ ;
wire \myidu/_0841_ ;
wire \myidu/_0842_ ;
wire \myidu/_0843_ ;
wire \myidu/_0844_ ;
wire \myidu/_0845_ ;
wire \myidu/_0846_ ;
wire \myidu/_0847_ ;
wire \myidu/_0848_ ;
wire \myidu/_0849_ ;
wire \myidu/_0850_ ;
wire \myidu/_0851_ ;
wire \myidu/_0852_ ;
wire \myidu/_0853_ ;
wire \myidu/_0854_ ;
wire \myidu/_0855_ ;
wire \myidu/_0856_ ;
wire \myidu/_0857_ ;
wire \myidu/_0858_ ;
wire \myidu/_0859_ ;
wire \myidu/_0860_ ;
wire \myidu/_0861_ ;
wire \myidu/_0862_ ;
wire \myidu/_0863_ ;
wire \myidu/_0864_ ;
wire \myidu/_0865_ ;
wire \myidu/_0866_ ;
wire \myidu/_0867_ ;
wire \myidu/_0868_ ;
wire \myidu/_0869_ ;
wire \myidu/_0870_ ;
wire \myidu/_0871_ ;
wire \myidu/_0872_ ;
wire \myidu/_0873_ ;
wire \myidu/_0874_ ;
wire \myidu/_0875_ ;
wire \myidu/_0876_ ;
wire \myidu/_0877_ ;
wire \myidu/_0878_ ;
wire \myidu/_0879_ ;
wire \myidu/_0880_ ;
wire \myidu/_0881_ ;
wire \myidu/_0882_ ;
wire \myidu/_0883_ ;
wire \myidu/_0884_ ;
wire \myidu/_0885_ ;
wire \myidu/_0886_ ;
wire \myidu/_0887_ ;
wire \myidu/_0888_ ;
wire \myidu/_0889_ ;
wire \myidu/_0890_ ;
wire \myidu/_0891_ ;
wire \myidu/_0892_ ;
wire \myidu/_0893_ ;
wire \myidu/_0894_ ;
wire \myidu/_0895_ ;
wire \myidu/_0896_ ;
wire \myidu/_0897_ ;
wire \myidu/_0898_ ;
wire \myidu/_0899_ ;
wire \myidu/_0900_ ;
wire \myidu/_0901_ ;
wire \myidu/_0902_ ;
wire \myidu/_0903_ ;
wire \myidu/_0904_ ;
wire \myidu/_0905_ ;
wire \myidu/_0906_ ;
wire \myidu/_0907_ ;
wire \myidu/_0908_ ;
wire \myidu/_0909_ ;
wire \myidu/_0910_ ;
wire \myidu/_0911_ ;
wire \myidu/_0912_ ;
wire \myidu/_0913_ ;
wire \myidu/_0914_ ;
wire \myidu/_0915_ ;
wire \myidu/_0916_ ;
wire \myidu/_0917_ ;
wire \myidu/_0918_ ;
wire \myidu/_0919_ ;
wire \myidu/_0920_ ;
wire \myidu/_0921_ ;
wire \myidu/_0922_ ;
wire \myidu/_0923_ ;
wire \myidu/_0924_ ;
wire \myidu/_0925_ ;
wire \myidu/_0926_ ;
wire \myidu/_0927_ ;
wire \myidu/_0928_ ;
wire \myidu/_0929_ ;
wire \myidu/_0930_ ;
wire \myidu/_0931_ ;
wire \myidu/_0932_ ;
wire \myidu/_0933_ ;
wire \myidu/_0934_ ;
wire \myidu/_0935_ ;
wire \myidu/_0936_ ;
wire \myidu/_0937_ ;
wire \myidu/_0938_ ;
wire \myidu/_0939_ ;
wire \myidu/_0940_ ;
wire \myidu/_0941_ ;
wire \myidu/_0942_ ;
wire \myidu/_0943_ ;
wire \myidu/_0944_ ;
wire \myidu/_0945_ ;
wire \myidu/_0946_ ;
wire \myidu/_0947_ ;
wire \myidu/_0948_ ;
wire \myidu/_0949_ ;
wire \myidu/_0950_ ;
wire \myidu/_0951_ ;
wire \myidu/_0952_ ;
wire \myidu/_0953_ ;
wire \myidu/_0954_ ;
wire \myidu/_0955_ ;
wire \myidu/_0956_ ;
wire \myidu/_0957_ ;
wire \myidu/_0958_ ;
wire \myidu/_0959_ ;
wire \myidu/_0960_ ;
wire \myidu/_0961_ ;
wire \myidu/_0962_ ;
wire \myidu/_0963_ ;
wire \myidu/_0964_ ;
wire \myidu/_0965_ ;
wire \myidu/_0966_ ;
wire \myidu/_0967_ ;
wire \myidu/_0968_ ;
wire \myidu/_0969_ ;
wire \myidu/_0970_ ;
wire \myidu/_0971_ ;
wire \myidu/_0972_ ;
wire \myidu/_0973_ ;
wire \myidu/_0974_ ;
wire \myidu/_0975_ ;
wire \myidu/_0976_ ;
wire \myidu/_0977_ ;
wire \myidu/_0978_ ;
wire \myidu/_0979_ ;
wire \myidu/_0980_ ;
wire \myidu/_0981_ ;
wire \myidu/_0982_ ;
wire \myidu/_0983_ ;
wire \myidu/_0984_ ;
wire \myidu/_0985_ ;
wire \myidu/_0986_ ;
wire \myidu/_0987_ ;
wire \myidu/_0988_ ;
wire \myidu/_0989_ ;
wire \myidu/_0990_ ;
wire \myidu/_0991_ ;
wire \myidu/_0992_ ;
wire \myidu/_0993_ ;
wire \myidu/_0994_ ;
wire \myidu/_0995_ ;
wire \myidu/_0996_ ;
wire \myidu/_0997_ ;
wire \myidu/_0998_ ;
wire \myidu/_0999_ ;
wire \myidu/_1000_ ;
wire \myidu/_1001_ ;
wire \myidu/_1002_ ;
wire \myidu/_1003_ ;
wire \myidu/_1004_ ;
wire \myidu/_1005_ ;
wire \myidu/_1006_ ;
wire \myidu/_1007_ ;
wire \myidu/_1008_ ;
wire \myifu/_0000_ ;
wire \myifu/_0001_ ;
wire \myifu/_0002_ ;
wire \myifu/_0003_ ;
wire \myifu/_0004_ ;
wire \myifu/_0005_ ;
wire \myifu/_0006_ ;
wire \myifu/_0007_ ;
wire \myifu/_0008_ ;
wire \myifu/_0009_ ;
wire \myifu/_0010_ ;
wire \myifu/_0011_ ;
wire \myifu/_0012_ ;
wire \myifu/_0013_ ;
wire \myifu/_0014_ ;
wire \myifu/_0015_ ;
wire \myifu/_0016_ ;
wire \myifu/_0017_ ;
wire \myifu/_0018_ ;
wire \myifu/_0019_ ;
wire \myifu/_0020_ ;
wire \myifu/_0021_ ;
wire \myifu/_0022_ ;
wire \myifu/_0023_ ;
wire \myifu/_0024_ ;
wire \myifu/_0025_ ;
wire \myifu/_0026_ ;
wire \myifu/_0027_ ;
wire \myifu/_0028_ ;
wire \myifu/_0029_ ;
wire \myifu/_0030_ ;
wire \myifu/_0031_ ;
wire \myifu/_0032_ ;
wire \myifu/_0033_ ;
wire \myifu/_0034_ ;
wire \myifu/_0035_ ;
wire \myifu/_0036_ ;
wire \myifu/_0037_ ;
wire \myifu/_0038_ ;
wire \myifu/_0039_ ;
wire \myifu/_0040_ ;
wire \myifu/_0041_ ;
wire \myifu/_0042_ ;
wire \myifu/_0043_ ;
wire \myifu/_0044_ ;
wire \myifu/_0045_ ;
wire \myifu/_0046_ ;
wire \myifu/_0047_ ;
wire \myifu/_0048_ ;
wire \myifu/_0049_ ;
wire \myifu/_0050_ ;
wire \myifu/_0051_ ;
wire \myifu/_0052_ ;
wire \myifu/_0053_ ;
wire \myifu/_0054_ ;
wire \myifu/_0055_ ;
wire \myifu/_0056_ ;
wire \myifu/_0057_ ;
wire \myifu/_0058_ ;
wire \myifu/_0059_ ;
wire \myifu/_0060_ ;
wire \myifu/_0061_ ;
wire \myifu/_0062_ ;
wire \myifu/_0063_ ;
wire \myifu/_0064_ ;
wire \myifu/_0065_ ;
wire \myifu/_0066_ ;
wire \myifu/_0067_ ;
wire \myifu/_0068_ ;
wire \myifu/_0069_ ;
wire \myifu/_0070_ ;
wire \myifu/_0071_ ;
wire \myifu/_0072_ ;
wire \myifu/_0073_ ;
wire \myifu/_0074_ ;
wire \myifu/_0075_ ;
wire \myifu/_0076_ ;
wire \myifu/_0077_ ;
wire \myifu/_0078_ ;
wire \myifu/_0079_ ;
wire \myifu/_0080_ ;
wire \myifu/_0081_ ;
wire \myifu/_0082_ ;
wire \myifu/_0083_ ;
wire \myifu/_0084_ ;
wire \myifu/_0085_ ;
wire \myifu/_0086_ ;
wire \myifu/_0087_ ;
wire \myifu/_0088_ ;
wire \myifu/_0089_ ;
wire \myifu/_0090_ ;
wire \myifu/_0091_ ;
wire \myifu/_0092_ ;
wire \myifu/_0093_ ;
wire \myifu/_0094_ ;
wire \myifu/_0095_ ;
wire \myifu/_0096_ ;
wire \myifu/_0097_ ;
wire \myifu/_0098_ ;
wire \myifu/_0099_ ;
wire \myifu/_0100_ ;
wire \myifu/_0101_ ;
wire \myifu/_0102_ ;
wire \myifu/_0103_ ;
wire \myifu/_0104_ ;
wire \myifu/_0105_ ;
wire \myifu/_0106_ ;
wire \myifu/_0107_ ;
wire \myifu/_0108_ ;
wire \myifu/_0109_ ;
wire \myifu/_0110_ ;
wire \myifu/_0111_ ;
wire \myifu/_0112_ ;
wire \myifu/_0113_ ;
wire \myifu/_0114_ ;
wire \myifu/_0115_ ;
wire \myifu/_0116_ ;
wire \myifu/_0117_ ;
wire \myifu/_0118_ ;
wire \myifu/_0119_ ;
wire \myifu/_0120_ ;
wire \myifu/_0121_ ;
wire \myifu/_0122_ ;
wire \myifu/_0123_ ;
wire \myifu/_0124_ ;
wire \myifu/_0125_ ;
wire \myifu/_0126_ ;
wire \myifu/_0127_ ;
wire \myifu/_0128_ ;
wire \myifu/_0129_ ;
wire \myifu/_0130_ ;
wire \myifu/_0131_ ;
wire \myifu/_0132_ ;
wire \myifu/_0133_ ;
wire \myifu/_0134_ ;
wire \myifu/_0135_ ;
wire \myifu/_0136_ ;
wire \myifu/_0137_ ;
wire \myifu/_0138_ ;
wire \myifu/_0139_ ;
wire \myifu/_0140_ ;
wire \myifu/_0141_ ;
wire \myifu/_0142_ ;
wire \myifu/_0143_ ;
wire \myifu/_0144_ ;
wire \myifu/_0145_ ;
wire \myifu/_0146_ ;
wire \myifu/_0147_ ;
wire \myifu/_0148_ ;
wire \myifu/_0149_ ;
wire \myifu/_0150_ ;
wire \myifu/_0151_ ;
wire \myifu/_0152_ ;
wire \myifu/_0153_ ;
wire \myifu/_0154_ ;
wire \myifu/_0155_ ;
wire \myifu/_0156_ ;
wire \myifu/_0157_ ;
wire \myifu/_0158_ ;
wire \myifu/_0159_ ;
wire \myifu/_0160_ ;
wire \myifu/_0161_ ;
wire \myifu/_0162_ ;
wire \myifu/_0163_ ;
wire \myifu/_0164_ ;
wire \myifu/_0165_ ;
wire \myifu/_0166_ ;
wire \myifu/_0167_ ;
wire \myifu/_0168_ ;
wire \myifu/_0169_ ;
wire \myifu/_0170_ ;
wire \myifu/_0171_ ;
wire \myifu/_0172_ ;
wire \myifu/_0173_ ;
wire \myifu/_0174_ ;
wire \myifu/_0175_ ;
wire \myifu/_0176_ ;
wire \myifu/_0177_ ;
wire \myifu/_0178_ ;
wire \myifu/_0179_ ;
wire \myifu/_0180_ ;
wire \myifu/_0181_ ;
wire \myifu/_0182_ ;
wire \myifu/_0183_ ;
wire \myifu/_0184_ ;
wire \myifu/_0185_ ;
wire \myifu/_0186_ ;
wire \myifu/_0187_ ;
wire \myifu/_0188_ ;
wire \myifu/_0189_ ;
wire \myifu/_0190_ ;
wire \myifu/_0191_ ;
wire \myifu/_0192_ ;
wire \myifu/_0193_ ;
wire \myifu/_0194_ ;
wire \myifu/_0195_ ;
wire \myifu/_0196_ ;
wire \myifu/_0197_ ;
wire \myifu/_0198_ ;
wire \myifu/_0199_ ;
wire \myifu/_0200_ ;
wire \myifu/_0201_ ;
wire \myifu/_0202_ ;
wire \myifu/_0203_ ;
wire \myifu/_0204_ ;
wire \myifu/_0205_ ;
wire \myifu/_0206_ ;
wire \myifu/_0207_ ;
wire \myifu/_0208_ ;
wire \myifu/_0209_ ;
wire \myifu/_0210_ ;
wire \myifu/_0211_ ;
wire \myifu/_0212_ ;
wire \myifu/_0213_ ;
wire \myifu/_0214_ ;
wire \myifu/_0215_ ;
wire \myifu/_0216_ ;
wire \myifu/_0217_ ;
wire \myifu/_0218_ ;
wire \myifu/_0219_ ;
wire \myifu/_0220_ ;
wire \myifu/_0221_ ;
wire \myifu/_0222_ ;
wire \myifu/_0223_ ;
wire \myifu/_0224_ ;
wire \myifu/_0225_ ;
wire \myifu/_0226_ ;
wire \myifu/_0227_ ;
wire \myifu/_0228_ ;
wire \myifu/_0229_ ;
wire \myifu/_0230_ ;
wire \myifu/_0231_ ;
wire \myifu/_0232_ ;
wire \myifu/_0233_ ;
wire \myifu/_0234_ ;
wire \myifu/_0235_ ;
wire \myifu/_0236_ ;
wire \myifu/_0237_ ;
wire \myifu/_0238_ ;
wire \myifu/_0239_ ;
wire \myifu/_0240_ ;
wire \myifu/_0241_ ;
wire \myifu/_0242_ ;
wire \myifu/_0243_ ;
wire \myifu/_0244_ ;
wire \myifu/_0245_ ;
wire \myifu/_0246_ ;
wire \myifu/_0247_ ;
wire \myifu/_0248_ ;
wire \myifu/_0249_ ;
wire \myifu/_0250_ ;
wire \myifu/_0251_ ;
wire \myifu/_0252_ ;
wire \myifu/_0253_ ;
wire \myifu/_0254_ ;
wire \myifu/_0255_ ;
wire \myifu/_0256_ ;
wire \myifu/_0257_ ;
wire \myifu/_0258_ ;
wire \myifu/_0259_ ;
wire \myifu/_0260_ ;
wire \myifu/_0261_ ;
wire \myifu/_0262_ ;
wire \myifu/_0263_ ;
wire \myifu/_0264_ ;
wire \myifu/_0265_ ;
wire \myifu/_0266_ ;
wire \myifu/_0267_ ;
wire \myifu/_0268_ ;
wire \myifu/_0269_ ;
wire \myifu/_0270_ ;
wire \myifu/_0271_ ;
wire \myifu/_0272_ ;
wire \myifu/_0273_ ;
wire \myifu/_0274_ ;
wire \myifu/_0275_ ;
wire \myifu/_0276_ ;
wire \myifu/_0277_ ;
wire \myifu/_0278_ ;
wire \myifu/_0279_ ;
wire \myifu/_0280_ ;
wire \myifu/_0281_ ;
wire \myifu/_0282_ ;
wire \myifu/_0283_ ;
wire \myifu/_0284_ ;
wire \myifu/_0285_ ;
wire \myifu/_0286_ ;
wire \myifu/_0287_ ;
wire \myifu/_0288_ ;
wire \myifu/_0289_ ;
wire \myifu/_0290_ ;
wire \myifu/_0291_ ;
wire \myifu/_0292_ ;
wire \myifu/_0293_ ;
wire \myifu/_0294_ ;
wire \myifu/_0295_ ;
wire \myifu/_0296_ ;
wire \myifu/_0297_ ;
wire \myifu/_0298_ ;
wire \myifu/_0299_ ;
wire \myifu/_0300_ ;
wire \myifu/_0301_ ;
wire \myifu/_0302_ ;
wire \myifu/_0303_ ;
wire \myifu/_0304_ ;
wire \myifu/_0305_ ;
wire \myifu/_0306_ ;
wire \myifu/_0307_ ;
wire \myifu/_0308_ ;
wire \myifu/_0309_ ;
wire \myifu/_0310_ ;
wire \myifu/_0311_ ;
wire \myifu/_0312_ ;
wire \myifu/_0313_ ;
wire \myifu/_0314_ ;
wire \myifu/_0315_ ;
wire \myifu/_0316_ ;
wire \myifu/_0317_ ;
wire \myifu/_0318_ ;
wire \myifu/_0319_ ;
wire \myifu/_0320_ ;
wire \myifu/_0321_ ;
wire \myifu/_0322_ ;
wire \myifu/_0323_ ;
wire \myifu/_0324_ ;
wire \myifu/_0325_ ;
wire \myifu/_0326_ ;
wire \myifu/_0327_ ;
wire \myifu/_0328_ ;
wire \myifu/_0329_ ;
wire \myifu/_0330_ ;
wire \myifu/_0331_ ;
wire \myifu/_0332_ ;
wire \myifu/_0333_ ;
wire \myifu/_0334_ ;
wire \myifu/_0335_ ;
wire \myifu/_0336_ ;
wire \myifu/_0337_ ;
wire \myifu/_0338_ ;
wire \myifu/_0339_ ;
wire \myifu/_0340_ ;
wire \myifu/_0341_ ;
wire \myifu/_0342_ ;
wire \myifu/_0343_ ;
wire \myifu/_0344_ ;
wire \myifu/_0345_ ;
wire \myifu/_0346_ ;
wire \myifu/_0347_ ;
wire \myifu/_0348_ ;
wire \myifu/_0349_ ;
wire \myifu/_0350_ ;
wire \myifu/_0351_ ;
wire \myifu/_0352_ ;
wire \myifu/_0353_ ;
wire \myifu/_0354_ ;
wire \myifu/_0355_ ;
wire \myifu/_0356_ ;
wire \myifu/_0357_ ;
wire \myifu/_0358_ ;
wire \myifu/_0359_ ;
wire \myifu/_0360_ ;
wire \myifu/_0361_ ;
wire \myifu/_0362_ ;
wire \myifu/_0363_ ;
wire \myifu/_0364_ ;
wire \myifu/_0365_ ;
wire \myifu/_0366_ ;
wire \myifu/_0367_ ;
wire \myifu/_0368_ ;
wire \myifu/_0369_ ;
wire \myifu/_0370_ ;
wire \myifu/_0371_ ;
wire \myifu/_0372_ ;
wire \myifu/_0373_ ;
wire \myifu/_0374_ ;
wire \myifu/_0375_ ;
wire \myifu/_0376_ ;
wire \myifu/_0377_ ;
wire \myifu/_0378_ ;
wire \myifu/_0379_ ;
wire \myifu/_0380_ ;
wire \myifu/_0381_ ;
wire \myifu/_0382_ ;
wire \myifu/_0383_ ;
wire \myifu/_0384_ ;
wire \myifu/_0385_ ;
wire \myifu/_0386_ ;
wire \myifu/_0387_ ;
wire \myifu/_0388_ ;
wire \myifu/_0389_ ;
wire \myifu/_0390_ ;
wire \myifu/_0391_ ;
wire \myifu/_0392_ ;
wire \myifu/_0393_ ;
wire \myifu/_0394_ ;
wire \myifu/_0395_ ;
wire \myifu/_0396_ ;
wire \myifu/_0397_ ;
wire \myifu/_0398_ ;
wire \myifu/_0399_ ;
wire \myifu/_0400_ ;
wire \myifu/_0401_ ;
wire \myifu/_0402_ ;
wire \myifu/_0403_ ;
wire \myifu/_0404_ ;
wire \myifu/_0405_ ;
wire \myifu/_0406_ ;
wire \myifu/_0407_ ;
wire \myifu/_0408_ ;
wire \myifu/_0409_ ;
wire \myifu/_0410_ ;
wire \myifu/_0411_ ;
wire \myifu/_0412_ ;
wire \myifu/_0413_ ;
wire \myifu/_0414_ ;
wire \myifu/_0415_ ;
wire \myifu/_0416_ ;
wire \myifu/_0417_ ;
wire \myifu/_0418_ ;
wire \myifu/_0419_ ;
wire \myifu/_0420_ ;
wire \myifu/_0421_ ;
wire \myifu/_0422_ ;
wire \myifu/_0423_ ;
wire \myifu/_0424_ ;
wire \myifu/_0425_ ;
wire \myifu/_0426_ ;
wire \myifu/_0427_ ;
wire \myifu/_0428_ ;
wire \myifu/_0429_ ;
wire \myifu/_0430_ ;
wire \myifu/_0431_ ;
wire \myifu/_0432_ ;
wire \myifu/_0433_ ;
wire \myifu/_0434_ ;
wire \myifu/_0435_ ;
wire \myifu/_0436_ ;
wire \myifu/_0437_ ;
wire \myifu/_0438_ ;
wire \myifu/_0439_ ;
wire \myifu/_0440_ ;
wire \myifu/_0441_ ;
wire \myifu/_0442_ ;
wire \myifu/_0443_ ;
wire \myifu/_0444_ ;
wire \myifu/_0445_ ;
wire \myifu/_0446_ ;
wire \myifu/_0447_ ;
wire \myifu/_0448_ ;
wire \myifu/_0449_ ;
wire \myifu/_0450_ ;
wire \myifu/_0451_ ;
wire \myifu/_0452_ ;
wire \myifu/_0453_ ;
wire \myifu/_0454_ ;
wire \myifu/_0455_ ;
wire \myifu/_0456_ ;
wire \myifu/_0457_ ;
wire \myifu/_0458_ ;
wire \myifu/_0459_ ;
wire \myifu/_0460_ ;
wire \myifu/_0461_ ;
wire \myifu/_0462_ ;
wire \myifu/_0463_ ;
wire \myifu/_0464_ ;
wire \myifu/_0465_ ;
wire \myifu/_0466_ ;
wire \myifu/_0467_ ;
wire \myifu/_0468_ ;
wire \myifu/_0469_ ;
wire \myifu/_0470_ ;
wire \myifu/_0471_ ;
wire \myifu/_0472_ ;
wire \myifu/_0473_ ;
wire \myifu/_0474_ ;
wire \myifu/_0475_ ;
wire \myifu/_0476_ ;
wire \myifu/_0477_ ;
wire \myifu/_0478_ ;
wire \myifu/_0479_ ;
wire \myifu/_0480_ ;
wire \myifu/_0481_ ;
wire \myifu/_0482_ ;
wire \myifu/_0483_ ;
wire \myifu/_0484_ ;
wire \myifu/_0485_ ;
wire \myifu/_0486_ ;
wire \myifu/_0487_ ;
wire \myifu/_0488_ ;
wire \myifu/_0489_ ;
wire \myifu/_0490_ ;
wire \myifu/_0491_ ;
wire \myifu/_0492_ ;
wire \myifu/_0493_ ;
wire \myifu/_0494_ ;
wire \myifu/_0495_ ;
wire \myifu/_0496_ ;
wire \myifu/_0497_ ;
wire \myifu/_0498_ ;
wire \myifu/_0499_ ;
wire \myifu/_0500_ ;
wire \myifu/_0501_ ;
wire \myifu/_0502_ ;
wire \myifu/_0503_ ;
wire \myifu/_0504_ ;
wire \myifu/_0505_ ;
wire \myifu/_0506_ ;
wire \myifu/_0507_ ;
wire \myifu/_0508_ ;
wire \myifu/_0509_ ;
wire \myifu/_0510_ ;
wire \myifu/_0511_ ;
wire \myifu/_0512_ ;
wire \myifu/_0513_ ;
wire \myifu/_0514_ ;
wire \myifu/_0515_ ;
wire \myifu/_0516_ ;
wire \myifu/_0517_ ;
wire \myifu/_0518_ ;
wire \myifu/_0519_ ;
wire \myifu/_0520_ ;
wire \myifu/_0521_ ;
wire \myifu/_0522_ ;
wire \myifu/_0523_ ;
wire \myifu/_0524_ ;
wire \myifu/_0525_ ;
wire \myifu/_0526_ ;
wire \myifu/_0527_ ;
wire \myifu/_0528_ ;
wire \myifu/_0529_ ;
wire \myifu/_0530_ ;
wire \myifu/_0531_ ;
wire \myifu/_0532_ ;
wire \myifu/_0533_ ;
wire \myifu/_0534_ ;
wire \myifu/_0535_ ;
wire \myifu/_0536_ ;
wire \myifu/_0537_ ;
wire \myifu/_0538_ ;
wire \myifu/_0539_ ;
wire \myifu/_0540_ ;
wire \myifu/_0541_ ;
wire \myifu/_0542_ ;
wire \myifu/_0543_ ;
wire \myifu/_0544_ ;
wire \myifu/_0545_ ;
wire \myifu/_0546_ ;
wire \myifu/_0547_ ;
wire \myifu/_0548_ ;
wire \myifu/_0549_ ;
wire \myifu/_0550_ ;
wire \myifu/_0551_ ;
wire \myifu/_0552_ ;
wire \myifu/_0553_ ;
wire \myifu/_0554_ ;
wire \myifu/_0555_ ;
wire \myifu/_0556_ ;
wire \myifu/_0557_ ;
wire \myifu/_0558_ ;
wire \myifu/_0559_ ;
wire \myifu/_0560_ ;
wire \myifu/_0561_ ;
wire \myifu/_0562_ ;
wire \myifu/_0563_ ;
wire \myifu/_0564_ ;
wire \myifu/_0565_ ;
wire \myifu/_0566_ ;
wire \myifu/_0567_ ;
wire \myifu/_0568_ ;
wire \myifu/_0569_ ;
wire \myifu/_0570_ ;
wire \myifu/_0571_ ;
wire \myifu/_0572_ ;
wire \myifu/_0573_ ;
wire \myifu/_0574_ ;
wire \myifu/_0575_ ;
wire \myifu/_0576_ ;
wire \myifu/_0577_ ;
wire \myifu/_0578_ ;
wire \myifu/_0579_ ;
wire \myifu/_0580_ ;
wire \myifu/_0581_ ;
wire \myifu/_0582_ ;
wire \myifu/_0583_ ;
wire \myifu/_0584_ ;
wire \myifu/_0585_ ;
wire \myifu/_0586_ ;
wire \myifu/_0587_ ;
wire \myifu/_0588_ ;
wire \myifu/_0589_ ;
wire \myifu/_0590_ ;
wire \myifu/_0591_ ;
wire \myifu/_0592_ ;
wire \myifu/_0593_ ;
wire \myifu/_0594_ ;
wire \myifu/_0595_ ;
wire \myifu/_0596_ ;
wire \myifu/_0597_ ;
wire \myifu/_0598_ ;
wire \myifu/_0599_ ;
wire \myifu/_0600_ ;
wire \myifu/_0601_ ;
wire \myifu/_0602_ ;
wire \myifu/_0603_ ;
wire \myifu/_0604_ ;
wire \myifu/_0605_ ;
wire \myifu/_0606_ ;
wire \myifu/_0607_ ;
wire \myifu/_0608_ ;
wire \myifu/_0609_ ;
wire \myifu/_0610_ ;
wire \myifu/_0611_ ;
wire \myifu/_0612_ ;
wire \myifu/_0613_ ;
wire \myifu/_0614_ ;
wire \myifu/_0615_ ;
wire \myifu/_0616_ ;
wire \myifu/_0617_ ;
wire \myifu/_0618_ ;
wire \myifu/_0619_ ;
wire \myifu/_0620_ ;
wire \myifu/_0621_ ;
wire \myifu/_0622_ ;
wire \myifu/_0623_ ;
wire \myifu/_0624_ ;
wire \myifu/_0625_ ;
wire \myifu/_0626_ ;
wire \myifu/_0627_ ;
wire \myifu/_0628_ ;
wire \myifu/_0629_ ;
wire \myifu/_0630_ ;
wire \myifu/_0631_ ;
wire \myifu/_0632_ ;
wire \myifu/_0633_ ;
wire \myifu/_0634_ ;
wire \myifu/_0635_ ;
wire \myifu/_0636_ ;
wire \myifu/_0637_ ;
wire \myifu/_0638_ ;
wire \myifu/_0639_ ;
wire \myifu/_0640_ ;
wire \myifu/_0641_ ;
wire \myifu/_0642_ ;
wire \myifu/_0643_ ;
wire \myifu/_0644_ ;
wire \myifu/_0645_ ;
wire \myifu/_0646_ ;
wire \myifu/_0647_ ;
wire \myifu/_0648_ ;
wire \myifu/_0649_ ;
wire \myifu/_0650_ ;
wire \myifu/_0651_ ;
wire \myifu/_0652_ ;
wire \myifu/_0653_ ;
wire \myifu/_0654_ ;
wire \myifu/_0655_ ;
wire \myifu/_0656_ ;
wire \myifu/_0657_ ;
wire \myifu/_0658_ ;
wire \myifu/_0659_ ;
wire \myifu/_0660_ ;
wire \myifu/_0661_ ;
wire \myifu/_0662_ ;
wire \myifu/_0663_ ;
wire \myifu/_0664_ ;
wire \myifu/_0665_ ;
wire \myifu/_0666_ ;
wire \myifu/_0667_ ;
wire \myifu/_0668_ ;
wire \myifu/_0669_ ;
wire \myifu/_0670_ ;
wire \myifu/_0671_ ;
wire \myifu/_0672_ ;
wire \myifu/_0673_ ;
wire \myifu/_0674_ ;
wire \myifu/_0675_ ;
wire \myifu/_0676_ ;
wire \myifu/_0677_ ;
wire \myifu/_0678_ ;
wire \myifu/_0679_ ;
wire \myifu/_0680_ ;
wire \myifu/_0681_ ;
wire \myifu/_0682_ ;
wire \myifu/_0683_ ;
wire \myifu/_0684_ ;
wire \myifu/_0685_ ;
wire \myifu/_0686_ ;
wire \myifu/_0687_ ;
wire \myifu/_0688_ ;
wire \myifu/_0689_ ;
wire \myifu/_0690_ ;
wire \myifu/_0691_ ;
wire \myifu/_0692_ ;
wire \myifu/_0693_ ;
wire \myifu/_0694_ ;
wire \myifu/_0695_ ;
wire \myifu/_0696_ ;
wire \myifu/_0697_ ;
wire \myifu/_0698_ ;
wire \myifu/_0699_ ;
wire \myifu/_0700_ ;
wire \myifu/_0701_ ;
wire \myifu/_0702_ ;
wire \myifu/_0703_ ;
wire \myifu/_0704_ ;
wire \myifu/_0705_ ;
wire \myifu/_0706_ ;
wire \myifu/_0707_ ;
wire \myifu/_0708_ ;
wire \myifu/_0709_ ;
wire \myifu/_0710_ ;
wire \myifu/_0711_ ;
wire \myifu/_0712_ ;
wire \myifu/_0713_ ;
wire \myifu/_0714_ ;
wire \myifu/_0715_ ;
wire \myifu/_0716_ ;
wire \myifu/_0717_ ;
wire \myifu/_0718_ ;
wire \myifu/_0719_ ;
wire \myifu/_0720_ ;
wire \myifu/_0721_ ;
wire \myifu/_0722_ ;
wire \myifu/_0723_ ;
wire \myifu/_0724_ ;
wire \myifu/_0725_ ;
wire \myifu/_0726_ ;
wire \myifu/_0727_ ;
wire \myifu/_0728_ ;
wire \myifu/_0729_ ;
wire \myifu/_0730_ ;
wire \myifu/_0731_ ;
wire \myifu/_0732_ ;
wire \myifu/_0733_ ;
wire \myifu/_0734_ ;
wire \myifu/_0735_ ;
wire \myifu/_0736_ ;
wire \myifu/_0737_ ;
wire \myifu/_0738_ ;
wire \myifu/_0739_ ;
wire \myifu/_0740_ ;
wire \myifu/_0741_ ;
wire \myifu/_0742_ ;
wire \myifu/_0743_ ;
wire \myifu/_0744_ ;
wire \myifu/_0745_ ;
wire \myifu/_0746_ ;
wire \myifu/_0747_ ;
wire \myifu/_0748_ ;
wire \myifu/_0749_ ;
wire \myifu/_0750_ ;
wire \myifu/_0751_ ;
wire \myifu/_0752_ ;
wire \myifu/_0753_ ;
wire \myifu/_0754_ ;
wire \myifu/_0755_ ;
wire \myifu/_0756_ ;
wire \myifu/_0757_ ;
wire \myifu/_0758_ ;
wire \myifu/_0759_ ;
wire \myifu/_0760_ ;
wire \myifu/_0761_ ;
wire \myifu/_0762_ ;
wire \myifu/_0763_ ;
wire \myifu/_0764_ ;
wire \myifu/_0765_ ;
wire \myifu/_0766_ ;
wire \myifu/_0767_ ;
wire \myifu/_0768_ ;
wire \myifu/_0769_ ;
wire \myifu/_0770_ ;
wire \myifu/_0771_ ;
wire \myifu/_0772_ ;
wire \myifu/_0773_ ;
wire \myifu/_0774_ ;
wire \myifu/_0775_ ;
wire \myifu/_0776_ ;
wire \myifu/_0777_ ;
wire \myifu/_0778_ ;
wire \myifu/_0779_ ;
wire \myifu/_0780_ ;
wire \myifu/_0781_ ;
wire \myifu/_0782_ ;
wire \myifu/_0783_ ;
wire \myifu/_0784_ ;
wire \myifu/_0785_ ;
wire \myifu/_0786_ ;
wire \myifu/_0787_ ;
wire \myifu/_0788_ ;
wire \myifu/_0789_ ;
wire \myifu/_0790_ ;
wire \myifu/_0791_ ;
wire \myifu/_0792_ ;
wire \myifu/_0793_ ;
wire \myifu/_0794_ ;
wire \myifu/_0795_ ;
wire \myifu/_0796_ ;
wire \myifu/_0797_ ;
wire \myifu/_0798_ ;
wire \myifu/_0799_ ;
wire \myifu/_0800_ ;
wire \myifu/_0801_ ;
wire \myifu/_0802_ ;
wire \myifu/_0803_ ;
wire \myifu/_0804_ ;
wire \myifu/_0805_ ;
wire \myifu/_0806_ ;
wire \myifu/_0807_ ;
wire \myifu/_0808_ ;
wire \myifu/_0809_ ;
wire \myifu/_0810_ ;
wire \myifu/_0811_ ;
wire \myifu/_0812_ ;
wire \myifu/_0813_ ;
wire \myifu/_0814_ ;
wire \myifu/_0815_ ;
wire \myifu/_0816_ ;
wire \myifu/_0817_ ;
wire \myifu/_0818_ ;
wire \myifu/_0819_ ;
wire \myifu/_0820_ ;
wire \myifu/_0821_ ;
wire \myifu/_0822_ ;
wire \myifu/_0823_ ;
wire \myifu/_0824_ ;
wire \myifu/_0825_ ;
wire \myifu/_0826_ ;
wire \myifu/_0827_ ;
wire \myifu/_0828_ ;
wire \myifu/_0829_ ;
wire \myifu/_0830_ ;
wire \myifu/_0831_ ;
wire \myifu/_0832_ ;
wire \myifu/_0833_ ;
wire \myifu/_0834_ ;
wire \myifu/_0835_ ;
wire \myifu/_0836_ ;
wire \myifu/_0837_ ;
wire \myifu/_0838_ ;
wire \myifu/_0839_ ;
wire \myifu/_0840_ ;
wire \myifu/_0841_ ;
wire \myifu/_0842_ ;
wire \myifu/_0843_ ;
wire \myifu/_0844_ ;
wire \myifu/_0845_ ;
wire \myifu/_0846_ ;
wire \myifu/_0847_ ;
wire \myifu/_0848_ ;
wire \myifu/_0849_ ;
wire \myifu/_0850_ ;
wire \myifu/_0851_ ;
wire \myifu/_0852_ ;
wire \myifu/_0853_ ;
wire \myifu/_0854_ ;
wire \myifu/_0855_ ;
wire \myifu/_0856_ ;
wire \myifu/_0857_ ;
wire \myifu/_0858_ ;
wire \myifu/_0859_ ;
wire \myifu/_0860_ ;
wire \myifu/_0861_ ;
wire \myifu/_0862_ ;
wire \myifu/_0863_ ;
wire \myifu/_0864_ ;
wire \myifu/_0865_ ;
wire \myifu/_0866_ ;
wire \myifu/_0867_ ;
wire \myifu/_0868_ ;
wire \myifu/_0869_ ;
wire \myifu/_0870_ ;
wire \myifu/_0871_ ;
wire \myifu/_0872_ ;
wire \myifu/_0873_ ;
wire \myifu/_0874_ ;
wire \myifu/_0875_ ;
wire \myifu/_0876_ ;
wire \myifu/_0877_ ;
wire \myifu/_0878_ ;
wire \myifu/_0879_ ;
wire \myifu/_0880_ ;
wire \myifu/_0881_ ;
wire \myifu/_0882_ ;
wire \myifu/_0883_ ;
wire \myifu/_0884_ ;
wire \myifu/_0885_ ;
wire \myifu/_0886_ ;
wire \myifu/_0887_ ;
wire \myifu/_0888_ ;
wire \myifu/_0889_ ;
wire \myifu/_0890_ ;
wire \myifu/_0891_ ;
wire \myifu/_0892_ ;
wire \myifu/_0893_ ;
wire \myifu/_0894_ ;
wire \myifu/_0895_ ;
wire \myifu/_0896_ ;
wire \myifu/_0897_ ;
wire \myifu/_0898_ ;
wire \myifu/_0899_ ;
wire \myifu/_0900_ ;
wire \myifu/_0901_ ;
wire \myifu/_0902_ ;
wire \myifu/_0903_ ;
wire \myifu/_0904_ ;
wire \myifu/_0905_ ;
wire \myifu/_0906_ ;
wire \myifu/_0907_ ;
wire \myifu/_0908_ ;
wire \myifu/_0909_ ;
wire \myifu/_0910_ ;
wire \myifu/_0911_ ;
wire \myifu/_0912_ ;
wire \myifu/_0913_ ;
wire \myifu/_0914_ ;
wire \myifu/_0915_ ;
wire \myifu/_0916_ ;
wire \myifu/_0917_ ;
wire \myifu/_0918_ ;
wire \myifu/_0919_ ;
wire \myifu/_0920_ ;
wire \myifu/_0921_ ;
wire \myifu/_0922_ ;
wire \myifu/_0923_ ;
wire \myifu/_0924_ ;
wire \myifu/_0925_ ;
wire \myifu/_0926_ ;
wire \myifu/_0927_ ;
wire \myifu/_0928_ ;
wire \myifu/_0929_ ;
wire \myifu/_0930_ ;
wire \myifu/_0931_ ;
wire \myifu/_0932_ ;
wire \myifu/_0933_ ;
wire \myifu/_0934_ ;
wire \myifu/_0935_ ;
wire \myifu/_0936_ ;
wire \myifu/_0937_ ;
wire \myifu/_0938_ ;
wire \myifu/_0939_ ;
wire \myifu/_0940_ ;
wire \myifu/_0941_ ;
wire \myifu/_0942_ ;
wire \myifu/_0943_ ;
wire \myifu/_0944_ ;
wire \myifu/_0945_ ;
wire \myifu/_0946_ ;
wire \myifu/_0947_ ;
wire \myifu/_0948_ ;
wire \myifu/_0949_ ;
wire \myifu/_0950_ ;
wire \myifu/_0951_ ;
wire \myifu/_0952_ ;
wire \myifu/_0953_ ;
wire \myifu/_0954_ ;
wire \myifu/_0955_ ;
wire \myifu/_0956_ ;
wire \myifu/_0957_ ;
wire \myifu/_0958_ ;
wire \myifu/_0959_ ;
wire \myifu/_0960_ ;
wire \myifu/_0961_ ;
wire \myifu/_0962_ ;
wire \myifu/_0963_ ;
wire \myifu/_0964_ ;
wire \myifu/_0965_ ;
wire \myifu/_0966_ ;
wire \myifu/_0967_ ;
wire \myifu/_0968_ ;
wire \myifu/_0969_ ;
wire \myifu/_0970_ ;
wire \myifu/_0971_ ;
wire \myifu/_0972_ ;
wire \myifu/_0973_ ;
wire \myifu/_0974_ ;
wire \myifu/_0975_ ;
wire \myifu/_0976_ ;
wire \myifu/_0977_ ;
wire \myifu/_0978_ ;
wire \myifu/_0979_ ;
wire \myifu/_0980_ ;
wire \myifu/_0981_ ;
wire \myifu/_0982_ ;
wire \myifu/_0983_ ;
wire \myifu/_0984_ ;
wire \myifu/_0985_ ;
wire \myifu/_0986_ ;
wire \myifu/_0987_ ;
wire \myifu/_0988_ ;
wire \myifu/_0989_ ;
wire \myifu/_0990_ ;
wire \myifu/_0991_ ;
wire \myifu/_0992_ ;
wire \myifu/_0993_ ;
wire \myifu/_0994_ ;
wire \myifu/_0995_ ;
wire \myifu/_0996_ ;
wire \myifu/_0997_ ;
wire \myifu/_0998_ ;
wire \myifu/_0999_ ;
wire \myifu/_1000_ ;
wire \myifu/_1001_ ;
wire \myifu/_1002_ ;
wire \myifu/_1003_ ;
wire \myifu/_1004_ ;
wire \myifu/_1005_ ;
wire \myifu/_1006_ ;
wire \myifu/_1007_ ;
wire \myifu/_1008_ ;
wire \myifu/_1009_ ;
wire \myifu/_1010_ ;
wire \myifu/_1011_ ;
wire \myifu/_1012_ ;
wire \myifu/_1013_ ;
wire \myifu/_1014_ ;
wire \myifu/_1015_ ;
wire \myifu/_1016_ ;
wire \myifu/_1017_ ;
wire \myifu/_1018_ ;
wire \myifu/_1019_ ;
wire \myifu/_1020_ ;
wire \myifu/_1021_ ;
wire \myifu/_1022_ ;
wire \myifu/_1023_ ;
wire \myifu/_1024_ ;
wire \myifu/_1025_ ;
wire \myifu/_1026_ ;
wire \myifu/_1027_ ;
wire \myifu/_1028_ ;
wire \myifu/_1029_ ;
wire \myifu/_1030_ ;
wire \myifu/_1031_ ;
wire \myifu/_1032_ ;
wire \myifu/_1033_ ;
wire \myifu/_1034_ ;
wire \myifu/_1035_ ;
wire \myifu/_1036_ ;
wire \myifu/_1037_ ;
wire \myifu/_1038_ ;
wire \myifu/_1039_ ;
wire \myifu/_1040_ ;
wire \myifu/_1041_ ;
wire \myifu/_1042_ ;
wire \myifu/_1043_ ;
wire \myifu/_1044_ ;
wire \myifu/_1045_ ;
wire \myifu/_1046_ ;
wire \myifu/_1047_ ;
wire \myifu/_1048_ ;
wire \myifu/_1049_ ;
wire \myifu/_1050_ ;
wire \myifu/_1051_ ;
wire \myifu/_1052_ ;
wire \myifu/_1053_ ;
wire \myifu/_1054_ ;
wire \myifu/_1055_ ;
wire \myifu/_1056_ ;
wire \myifu/_1057_ ;
wire \myifu/_1058_ ;
wire \myifu/_1059_ ;
wire \myifu/_1060_ ;
wire \myifu/_1061_ ;
wire \myifu/_1062_ ;
wire \myifu/_1063_ ;
wire \myifu/_1064_ ;
wire \myifu/_1065_ ;
wire \myifu/_1066_ ;
wire \myifu/_1067_ ;
wire \myifu/_1068_ ;
wire \myifu/_1069_ ;
wire \myifu/_1070_ ;
wire \myifu/_1071_ ;
wire \myifu/_1072_ ;
wire \myifu/_1073_ ;
wire \myifu/_1074_ ;
wire \myifu/_1075_ ;
wire \myifu/_1076_ ;
wire \myifu/_1077_ ;
wire \myifu/_1078_ ;
wire \myifu/_1079_ ;
wire \myifu/_1080_ ;
wire \myifu/_1081_ ;
wire \myifu/_1082_ ;
wire \myifu/_1083_ ;
wire \myifu/_1084_ ;
wire \myifu/_1085_ ;
wire \myifu/_1086_ ;
wire \myifu/_1087_ ;
wire \myifu/_1088_ ;
wire \myifu/_1089_ ;
wire \myifu/_1090_ ;
wire \myifu/_1091_ ;
wire \myifu/_1092_ ;
wire \myifu/_1093_ ;
wire \myifu/_1094_ ;
wire \myifu/_1095_ ;
wire \myifu/_1096_ ;
wire \myifu/_1097_ ;
wire \myifu/pred_jump ;
wire \myifu/valid_in ;
wire \myifu/valid_out ;
wire \myifu/myicache/_0000_ ;
wire \myifu/myicache/_0001_ ;
wire \myifu/myicache/_0002_ ;
wire \myifu/myicache/_0003_ ;
wire \myifu/myicache/_0004_ ;
wire \myifu/myicache/_0005_ ;
wire \myifu/myicache/_0006_ ;
wire \myifu/myicache/_0007_ ;
wire \myifu/myicache/_0008_ ;
wire \myifu/myicache/_0009_ ;
wire \myifu/myicache/_0010_ ;
wire \myifu/myicache/_0011_ ;
wire \myifu/myicache/_0012_ ;
wire \myifu/myicache/_0013_ ;
wire \myifu/myicache/_0014_ ;
wire \myifu/myicache/_0015_ ;
wire \myifu/myicache/_0016_ ;
wire \myifu/myicache/_0017_ ;
wire \myifu/myicache/_0018_ ;
wire \myifu/myicache/_0019_ ;
wire \myifu/myicache/_0020_ ;
wire \myifu/myicache/_0021_ ;
wire \myifu/myicache/_0022_ ;
wire \myifu/myicache/_0023_ ;
wire \myifu/myicache/_0024_ ;
wire \myifu/myicache/_0025_ ;
wire \myifu/myicache/_0026_ ;
wire \myifu/myicache/_0027_ ;
wire \myifu/myicache/_0028_ ;
wire \myifu/myicache/_0029_ ;
wire \myifu/myicache/_0030_ ;
wire \myifu/myicache/_0031_ ;
wire \myifu/myicache/_0032_ ;
wire \myifu/myicache/_0033_ ;
wire \myifu/myicache/_0034_ ;
wire \myifu/myicache/_0035_ ;
wire \myifu/myicache/_0036_ ;
wire \myifu/myicache/_0037_ ;
wire \myifu/myicache/_0038_ ;
wire \myifu/myicache/_0039_ ;
wire \myifu/myicache/_0040_ ;
wire \myifu/myicache/_0041_ ;
wire \myifu/myicache/_0042_ ;
wire \myifu/myicache/_0043_ ;
wire \myifu/myicache/_0044_ ;
wire \myifu/myicache/_0045_ ;
wire \myifu/myicache/_0046_ ;
wire \myifu/myicache/_0047_ ;
wire \myifu/myicache/_0048_ ;
wire \myifu/myicache/_0049_ ;
wire \myifu/myicache/_0050_ ;
wire \myifu/myicache/_0051_ ;
wire \myifu/myicache/_0052_ ;
wire \myifu/myicache/_0053_ ;
wire \myifu/myicache/_0054_ ;
wire \myifu/myicache/_0055_ ;
wire \myifu/myicache/_0056_ ;
wire \myifu/myicache/_0057_ ;
wire \myifu/myicache/_0058_ ;
wire \myifu/myicache/_0059_ ;
wire \myifu/myicache/_0060_ ;
wire \myifu/myicache/_0061_ ;
wire \myifu/myicache/_0062_ ;
wire \myifu/myicache/_0063_ ;
wire \myifu/myicache/_0064_ ;
wire \myifu/myicache/_0065_ ;
wire \myifu/myicache/_0066_ ;
wire \myifu/myicache/_0067_ ;
wire \myifu/myicache/_0068_ ;
wire \myifu/myicache/_0069_ ;
wire \myifu/myicache/_0070_ ;
wire \myifu/myicache/_0071_ ;
wire \myifu/myicache/_0072_ ;
wire \myifu/myicache/_0073_ ;
wire \myifu/myicache/_0074_ ;
wire \myifu/myicache/_0075_ ;
wire \myifu/myicache/_0076_ ;
wire \myifu/myicache/_0077_ ;
wire \myifu/myicache/_0078_ ;
wire \myifu/myicache/_0079_ ;
wire \myifu/myicache/_0080_ ;
wire \myifu/myicache/_0081_ ;
wire \myifu/myicache/_0082_ ;
wire \myifu/myicache/_0083_ ;
wire \myifu/myicache/_0084_ ;
wire \myifu/myicache/_0085_ ;
wire \myifu/myicache/_0086_ ;
wire \myifu/myicache/_0087_ ;
wire \myifu/myicache/_0088_ ;
wire \myifu/myicache/_0089_ ;
wire \myifu/myicache/_0090_ ;
wire \myifu/myicache/_0091_ ;
wire \myifu/myicache/_0092_ ;
wire \myifu/myicache/_0093_ ;
wire \myifu/myicache/_0094_ ;
wire \myifu/myicache/_0095_ ;
wire \myifu/myicache/_0096_ ;
wire \myifu/myicache/_0097_ ;
wire \myifu/myicache/_0098_ ;
wire \myifu/myicache/_0099_ ;
wire \myifu/myicache/_0100_ ;
wire \myifu/myicache/_0101_ ;
wire \myifu/myicache/_0102_ ;
wire \myifu/myicache/_0103_ ;
wire \myifu/myicache/_0104_ ;
wire \myifu/myicache/_0105_ ;
wire \myifu/myicache/_0106_ ;
wire \myifu/myicache/_0107_ ;
wire \myifu/myicache/_0108_ ;
wire \myifu/myicache/_0109_ ;
wire \myifu/myicache/_0110_ ;
wire \myifu/myicache/_0111_ ;
wire \myifu/myicache/_0112_ ;
wire \myifu/myicache/_0113_ ;
wire \myifu/myicache/_0114_ ;
wire \myifu/myicache/_0115_ ;
wire \myifu/myicache/_0116_ ;
wire \myifu/myicache/_0117_ ;
wire \myifu/myicache/_0118_ ;
wire \myifu/myicache/_0119_ ;
wire \myifu/myicache/_0120_ ;
wire \myifu/myicache/_0121_ ;
wire \myifu/myicache/_0122_ ;
wire \myifu/myicache/_0123_ ;
wire \myifu/myicache/_0124_ ;
wire \myifu/myicache/_0125_ ;
wire \myifu/myicache/_0126_ ;
wire \myifu/myicache/_0127_ ;
wire \myifu/myicache/_0128_ ;
wire \myifu/myicache/_0129_ ;
wire \myifu/myicache/_0130_ ;
wire \myifu/myicache/_0131_ ;
wire \myifu/myicache/_0132_ ;
wire \myifu/myicache/_0133_ ;
wire \myifu/myicache/_0134_ ;
wire \myifu/myicache/_0135_ ;
wire \myifu/myicache/_0136_ ;
wire \myifu/myicache/_0137_ ;
wire \myifu/myicache/_0138_ ;
wire \myifu/myicache/_0139_ ;
wire \myifu/myicache/_0140_ ;
wire \myifu/myicache/_0141_ ;
wire \myifu/myicache/_0142_ ;
wire \myifu/myicache/_0143_ ;
wire \myifu/myicache/_0144_ ;
wire \myifu/myicache/_0145_ ;
wire \myifu/myicache/_0146_ ;
wire \myifu/myicache/_0147_ ;
wire \myifu/myicache/_0148_ ;
wire \myifu/myicache/_0149_ ;
wire \myifu/myicache/_0150_ ;
wire \myifu/myicache/_0151_ ;
wire \myifu/myicache/_0152_ ;
wire \myifu/myicache/_0153_ ;
wire \myifu/myicache/_0154_ ;
wire \myifu/myicache/_0155_ ;
wire \myifu/myicache/_0156_ ;
wire \myifu/myicache/_0157_ ;
wire \myifu/myicache/_0158_ ;
wire \myifu/myicache/_0159_ ;
wire \myifu/myicache/_0160_ ;
wire \myifu/myicache/_0161_ ;
wire \myifu/myicache/_0162_ ;
wire \myifu/myicache/_0163_ ;
wire \myifu/myicache/_0164_ ;
wire \myifu/myicache/_0165_ ;
wire \myifu/myicache/_0166_ ;
wire \myifu/myicache/_0167_ ;
wire \myifu/myicache/_0168_ ;
wire \myifu/myicache/_0169_ ;
wire \myifu/myicache/_0170_ ;
wire \myifu/myicache/_0171_ ;
wire \myifu/myicache/_0172_ ;
wire \myifu/myicache/_0173_ ;
wire \myifu/myicache/_0174_ ;
wire \myifu/myicache/_0175_ ;
wire \myifu/myicache/_0176_ ;
wire \myifu/myicache/_0177_ ;
wire \myifu/myicache/_0178_ ;
wire \myifu/myicache/_0179_ ;
wire \myifu/myicache/_0180_ ;
wire \myifu/myicache/_0181_ ;
wire \myifu/myicache/_0182_ ;
wire \myifu/myicache/_0183_ ;
wire \myifu/myicache/_0184_ ;
wire \myifu/myicache/_0185_ ;
wire \myifu/myicache/_0186_ ;
wire \myifu/myicache/_0187_ ;
wire \myifu/myicache/_0188_ ;
wire \myifu/myicache/_0189_ ;
wire \myifu/myicache/_0190_ ;
wire \myifu/myicache/_0191_ ;
wire \myifu/myicache/_0192_ ;
wire \myifu/myicache/_0193_ ;
wire \myifu/myicache/_0194_ ;
wire \myifu/myicache/_0195_ ;
wire \myifu/myicache/_0196_ ;
wire \myifu/myicache/_0197_ ;
wire \myifu/myicache/_0198_ ;
wire \myifu/myicache/_0199_ ;
wire \myifu/myicache/_0200_ ;
wire \myifu/myicache/_0201_ ;
wire \myifu/myicache/_0202_ ;
wire \myifu/myicache/_0203_ ;
wire \myifu/myicache/_0204_ ;
wire \myifu/myicache/_0205_ ;
wire \myifu/myicache/_0206_ ;
wire \myifu/myicache/_0207_ ;
wire \myifu/myicache/_0208_ ;
wire \myifu/myicache/_0209_ ;
wire \myifu/myicache/_0210_ ;
wire \myifu/myicache/_0211_ ;
wire \myifu/myicache/_0212_ ;
wire \myifu/myicache/_0213_ ;
wire \myifu/myicache/_0214_ ;
wire \myifu/myicache/_0215_ ;
wire \myifu/myicache/_0216_ ;
wire \myifu/myicache/_0217_ ;
wire \myifu/myicache/_0218_ ;
wire \myifu/myicache/_0219_ ;
wire \myifu/myicache/_0220_ ;
wire \myifu/myicache/_0221_ ;
wire \myifu/myicache/_0222_ ;
wire \myifu/myicache/_0223_ ;
wire \myifu/myicache/_0224_ ;
wire \myifu/myicache/_0225_ ;
wire \myifu/myicache/_0226_ ;
wire \myifu/myicache/_0227_ ;
wire \myifu/myicache/_0228_ ;
wire \myifu/myicache/_0229_ ;
wire \myifu/myicache/_0230_ ;
wire \myifu/myicache/_0231_ ;
wire \myifu/myicache/_0232_ ;
wire \myifu/myicache/_0233_ ;
wire \myifu/myicache/_0234_ ;
wire \myifu/myicache/_0235_ ;
wire \myifu/myicache/_0236_ ;
wire \myifu/myicache/_0237_ ;
wire \myifu/myicache/_0238_ ;
wire \myifu/myicache/_0239_ ;
wire \myifu/myicache/_0240_ ;
wire \myifu/myicache/_0241_ ;
wire \myifu/myicache/_0242_ ;
wire \myifu/myicache/_0243_ ;
wire \myifu/myicache/_0244_ ;
wire \myifu/myicache/_0245_ ;
wire \myifu/myicache/_0246_ ;
wire \myifu/myicache/_0247_ ;
wire \myifu/myicache/_0248_ ;
wire \myifu/myicache/_0249_ ;
wire \myifu/myicache/_0250_ ;
wire \myifu/myicache/_0251_ ;
wire \myifu/myicache/_0252_ ;
wire \myifu/myicache/_0253_ ;
wire \myifu/myicache/_0254_ ;
wire \myifu/myicache/_0255_ ;
wire \myifu/myicache/_0256_ ;
wire \myifu/myicache/_0257_ ;
wire \myifu/myicache/_0258_ ;
wire \myifu/myicache/_0259_ ;
wire \myifu/myicache/_0260_ ;
wire \myifu/myicache/_0261_ ;
wire \myifu/myicache/_0262_ ;
wire \myifu/myicache/_0263_ ;
wire \myifu/myicache/_0264_ ;
wire \myifu/myicache/_0265_ ;
wire \myifu/myicache/_0266_ ;
wire \myifu/myicache/_0267_ ;
wire \myifu/myicache/_0268_ ;
wire \myifu/myicache/_0269_ ;
wire \myifu/myicache/_0270_ ;
wire \myifu/myicache/_0271_ ;
wire \myifu/myicache/_0272_ ;
wire \myifu/myicache/_0273_ ;
wire \myifu/myicache/_0274_ ;
wire \myifu/myicache/_0275_ ;
wire \myifu/myicache/_0276_ ;
wire \myifu/myicache/_0277_ ;
wire \myifu/myicache/_0278_ ;
wire \myifu/myicache/_0279_ ;
wire \myifu/myicache/_0280_ ;
wire \myifu/myicache/_0281_ ;
wire \myifu/myicache/_0282_ ;
wire \myifu/myicache/_0283_ ;
wire \myifu/myicache/_0284_ ;
wire \myifu/myicache/_0285_ ;
wire \myifu/myicache/_0286_ ;
wire \myifu/myicache/_0287_ ;
wire \myifu/myicache/_0288_ ;
wire \myifu/myicache/_0289_ ;
wire \myifu/myicache/_0290_ ;
wire \myifu/myicache/_0291_ ;
wire \myifu/myicache/_0292_ ;
wire \myifu/myicache/_0293_ ;
wire \myifu/myicache/_0294_ ;
wire \myifu/myicache/_0295_ ;
wire \myifu/myicache/_0296_ ;
wire \myifu/myicache/_0297_ ;
wire \myifu/myicache/_0298_ ;
wire \myifu/myicache/_0299_ ;
wire \myifu/myicache/_0300_ ;
wire \myifu/myicache/_0301_ ;
wire \myifu/myicache/_0302_ ;
wire \myifu/myicache/_0303_ ;
wire \myifu/myicache/_0304_ ;
wire \myifu/myicache/_0305_ ;
wire \myifu/myicache/_0306_ ;
wire \myifu/myicache/_0307_ ;
wire \myifu/myicache/_0308_ ;
wire \myifu/myicache/_0309_ ;
wire \myifu/myicache/_0310_ ;
wire \myifu/myicache/_0311_ ;
wire \myifu/myicache/_0312_ ;
wire \myifu/myicache/_0313_ ;
wire \myifu/myicache/_0314_ ;
wire \myifu/myicache/_0315_ ;
wire \myifu/myicache/_0316_ ;
wire \myifu/myicache/_0317_ ;
wire \myifu/myicache/_0318_ ;
wire \myifu/myicache/_0319_ ;
wire \myifu/myicache/_0320_ ;
wire \myifu/myicache/_0321_ ;
wire \myifu/myicache/_0322_ ;
wire \myifu/myicache/_0323_ ;
wire \myifu/myicache/_0324_ ;
wire \myifu/myicache/_0325_ ;
wire \myifu/myicache/_0326_ ;
wire \myifu/myicache/_0327_ ;
wire \myifu/myicache/_0328_ ;
wire \myifu/myicache/_0329_ ;
wire \myifu/myicache/_0330_ ;
wire \myifu/myicache/_0331_ ;
wire \myifu/myicache/_0332_ ;
wire \myifu/myicache/_0333_ ;
wire \myifu/myicache/_0334_ ;
wire \myifu/myicache/_0335_ ;
wire \myifu/myicache/_0336_ ;
wire \myifu/myicache/_0337_ ;
wire \myifu/myicache/_0338_ ;
wire \myifu/myicache/_0339_ ;
wire \myifu/myicache/_0340_ ;
wire \myifu/myicache/_0341_ ;
wire \myifu/myicache/_0342_ ;
wire \myifu/myicache/_0343_ ;
wire \myifu/myicache/_0344_ ;
wire \myifu/myicache/_0345_ ;
wire \myifu/myicache/_0346_ ;
wire \myifu/myicache/_0347_ ;
wire \myifu/myicache/_0348_ ;
wire \myifu/myicache/_0349_ ;
wire \myifu/myicache/_0350_ ;
wire \myifu/myicache/_0351_ ;
wire \myifu/myicache/_0352_ ;
wire \myifu/myicache/_0353_ ;
wire \myifu/myicache/_0354_ ;
wire \myifu/myicache/_0355_ ;
wire \myifu/myicache/_0356_ ;
wire \myifu/myicache/_0357_ ;
wire \myifu/myicache/_0358_ ;
wire \myifu/myicache/_0359_ ;
wire \myifu/myicache/_0360_ ;
wire \myifu/myicache/_0361_ ;
wire \myifu/myicache/_0362_ ;
wire \myifu/myicache/_0363_ ;
wire \myifu/myicache/_0364_ ;
wire \myifu/myicache/_0365_ ;
wire \myifu/myicache/_0366_ ;
wire \myifu/myicache/_0367_ ;
wire \myifu/myicache/_0368_ ;
wire \myifu/myicache/_0369_ ;
wire \myifu/myicache/_0370_ ;
wire \myifu/myicache/_0371_ ;
wire \myifu/myicache/_0372_ ;
wire \myifu/myicache/_0373_ ;
wire \myifu/myicache/_0374_ ;
wire \myifu/myicache/_0375_ ;
wire \myifu/myicache/_0376_ ;
wire \myifu/myicache/_0377_ ;
wire \myifu/myicache/_0378_ ;
wire \myifu/myicache/_0379_ ;
wire \myifu/myicache/_0380_ ;
wire \myifu/myicache/_0381_ ;
wire \myifu/myicache/_0382_ ;
wire \myifu/myicache/_0383_ ;
wire \myifu/myicache/_0384_ ;
wire \myifu/myicache/_0385_ ;
wire \myifu/myicache/_0386_ ;
wire \myifu/myicache/_0387_ ;
wire \myifu/myicache/_0388_ ;
wire \myifu/myicache/_0389_ ;
wire \myifu/myicache/_0390_ ;
wire \myifu/myicache/_0391_ ;
wire \myifu/myicache/_0392_ ;
wire \myifu/myicache/_0393_ ;
wire \myifu/myicache/_0394_ ;
wire \myifu/myicache/_0395_ ;
wire \myifu/myicache/_0396_ ;
wire \myifu/myicache/_0397_ ;
wire \myifu/myicache/_0398_ ;
wire \myifu/myicache/_0399_ ;
wire \myifu/myicache/_0400_ ;
wire \myifu/myicache/_0401_ ;
wire \myifu/myicache/_0402_ ;
wire \myifu/myicache/_0403_ ;
wire \myifu/myicache/_0404_ ;
wire \myifu/myicache/_0405_ ;
wire \myifu/myicache/_0406_ ;
wire \myifu/myicache/_0407_ ;
wire \myifu/myicache/_0408_ ;
wire \myifu/myicache/_0409_ ;
wire \myifu/myicache/_0410_ ;
wire \myifu/myicache/_0411_ ;
wire \myifu/myicache/_0412_ ;
wire \myifu/myicache/_0413_ ;
wire \myifu/myicache/_0414_ ;
wire \myifu/myicache/_0415_ ;
wire \myifu/myicache/_0416_ ;
wire \myifu/myicache/_0417_ ;
wire \myifu/myicache/_0418_ ;
wire \myifu/myicache/_0419_ ;
wire \myifu/myicache/_0420_ ;
wire \myifu/myicache/_0421_ ;
wire \myifu/myicache/_0422_ ;
wire \myifu/myicache/_0423_ ;
wire \myifu/myicache/_0424_ ;
wire \myifu/myicache/_0425_ ;
wire \myifu/myicache/_0426_ ;
wire \myifu/myicache/_0427_ ;
wire \myifu/myicache/_0428_ ;
wire \myifu/myicache/_0429_ ;
wire \myifu/myicache/_0430_ ;
wire \myifu/myicache/_0431_ ;
wire \myifu/myicache/_0432_ ;
wire \myifu/myicache/_0433_ ;
wire \myifu/myicache/_0434_ ;
wire \myifu/myicache/_0435_ ;
wire \myifu/myicache/_0436_ ;
wire \myifu/myicache/_0437_ ;
wire \myifu/myicache/_0438_ ;
wire \myifu/myicache/_0439_ ;
wire \myifu/myicache/_0440_ ;
wire \myifu/myicache/_0441_ ;
wire \myifu/myicache/_0442_ ;
wire \myifu/myicache/_0443_ ;
wire \myifu/myicache/_0444_ ;
wire \myifu/myicache/_0445_ ;
wire \myifu/myicache/_0446_ ;
wire \myifu/myicache/_0447_ ;
wire \myifu/myicache/_0448_ ;
wire \myifu/myicache/_0449_ ;
wire \myifu/myicache/_0450_ ;
wire \myifu/myicache/_0451_ ;
wire \myifu/myicache/_0452_ ;
wire \myifu/myicache/_0453_ ;
wire \myifu/myicache/_0454_ ;
wire \myifu/myicache/_0455_ ;
wire \myifu/myicache/_0456_ ;
wire \myifu/myicache/_0457_ ;
wire \myifu/myicache/_0458_ ;
wire \myifu/myicache/_0459_ ;
wire \myifu/myicache/_0460_ ;
wire \myifu/myicache/_0461_ ;
wire \myifu/myicache/_0462_ ;
wire \myifu/myicache/_0463_ ;
wire \myifu/myicache/_0464_ ;
wire \myifu/myicache/_0465_ ;
wire \myifu/myicache/_0466_ ;
wire \myifu/myicache/_0467_ ;
wire \myifu/myicache/_0468_ ;
wire \myifu/myicache/_0469_ ;
wire \myifu/myicache/_0470_ ;
wire \myifu/myicache/_0471_ ;
wire \myifu/myicache/_0472_ ;
wire \myifu/myicache/_0473_ ;
wire \myifu/myicache/_0474_ ;
wire \myifu/myicache/_0475_ ;
wire \myifu/myicache/_0476_ ;
wire \myifu/myicache/_0477_ ;
wire \myifu/myicache/_0478_ ;
wire \myifu/myicache/_0479_ ;
wire \myifu/myicache/_0480_ ;
wire \myifu/myicache/_0481_ ;
wire \myifu/myicache/_0482_ ;
wire \myifu/myicache/_0483_ ;
wire \myifu/myicache/_0484_ ;
wire \myifu/myicache/_0485_ ;
wire \myifu/myicache/_0486_ ;
wire \myifu/myicache/_0487_ ;
wire \myifu/myicache/_0488_ ;
wire \myifu/myicache/_0489_ ;
wire \myifu/myicache/_0490_ ;
wire \myifu/myicache/_0491_ ;
wire \myifu/myicache/_0492_ ;
wire \myifu/myicache/_0493_ ;
wire \myifu/myicache/_0494_ ;
wire \myifu/myicache/_0495_ ;
wire \myifu/myicache/_0496_ ;
wire \myifu/myicache/_0497_ ;
wire \myifu/myicache/_0498_ ;
wire \myifu/myicache/_0499_ ;
wire \myifu/myicache/_0500_ ;
wire \myifu/myicache/_0501_ ;
wire \myifu/myicache/_0502_ ;
wire \myifu/myicache/_0503_ ;
wire \myifu/myicache/_0504_ ;
wire \myifu/myicache/_0505_ ;
wire \myifu/myicache/_0506_ ;
wire \myifu/myicache/_0507_ ;
wire \myifu/myicache/_0508_ ;
wire \myifu/myicache/_0509_ ;
wire \myifu/myicache/_0510_ ;
wire \myifu/myicache/_0511_ ;
wire \myifu/myicache/_0512_ ;
wire \myifu/myicache/_0513_ ;
wire \myifu/myicache/_0514_ ;
wire \myifu/myicache/_0515_ ;
wire \myifu/myicache/_0516_ ;
wire \myifu/myicache/_0517_ ;
wire \myifu/myicache/_0518_ ;
wire \myifu/myicache/_0519_ ;
wire \myifu/myicache/_0520_ ;
wire \myifu/myicache/_0521_ ;
wire \myifu/myicache/_0522_ ;
wire \myifu/myicache/_0523_ ;
wire \myifu/myicache/_0524_ ;
wire \myifu/myicache/_0525_ ;
wire \myifu/myicache/_0526_ ;
wire \myifu/myicache/_0527_ ;
wire \myifu/myicache/_0528_ ;
wire \myifu/myicache/_0529_ ;
wire \myifu/myicache/_0530_ ;
wire \myifu/myicache/_0531_ ;
wire \myifu/myicache/_0532_ ;
wire \myifu/myicache/_0533_ ;
wire \myifu/myicache/_0534_ ;
wire \myifu/myicache/_0535_ ;
wire \myifu/myicache/_0536_ ;
wire \myifu/myicache/_0537_ ;
wire \myifu/myicache/_0538_ ;
wire \myifu/myicache/_0539_ ;
wire \myifu/myicache/_0540_ ;
wire \myifu/myicache/_0541_ ;
wire \myifu/myicache/_0542_ ;
wire \myifu/myicache/_0543_ ;
wire \myifu/myicache/_0544_ ;
wire \myifu/myicache/_0545_ ;
wire \myifu/myicache/_0546_ ;
wire \myifu/myicache/_0547_ ;
wire \myifu/myicache/_0548_ ;
wire \myifu/myicache/_0549_ ;
wire \myifu/myicache/_0550_ ;
wire \myifu/myicache/_0551_ ;
wire \myifu/myicache/_0552_ ;
wire \myifu/myicache/_0553_ ;
wire \myifu/myicache/_0554_ ;
wire \myifu/myicache/_0555_ ;
wire \myifu/myicache/_0556_ ;
wire \myifu/myicache/_0557_ ;
wire \myifu/myicache/_0558_ ;
wire \myifu/myicache/_0559_ ;
wire \myifu/myicache/_0560_ ;
wire \myifu/myicache/_0561_ ;
wire \myifu/myicache/_0562_ ;
wire \myifu/myicache/_0563_ ;
wire \myifu/myicache/_0564_ ;
wire \myifu/myicache/_0565_ ;
wire \myifu/myicache/_0566_ ;
wire \myifu/myicache/_0567_ ;
wire \myifu/myicache/_0568_ ;
wire \myifu/myicache/_0569_ ;
wire \myifu/myicache/_0570_ ;
wire \myifu/myicache/_0571_ ;
wire \myifu/myicache/_0572_ ;
wire \myifu/myicache/_0573_ ;
wire \myifu/myicache/_0574_ ;
wire \myifu/myicache/_0575_ ;
wire \myifu/myicache/_0576_ ;
wire \myifu/myicache/_0577_ ;
wire \myifu/myicache/_0578_ ;
wire \myifu/myicache/_0579_ ;
wire \myifu/myicache/_0580_ ;
wire \myifu/myicache/_0581_ ;
wire \myifu/myicache/_0582_ ;
wire \myifu/myicache/_0583_ ;
wire \myifu/myicache/_0584_ ;
wire \myifu/myicache/_0585_ ;
wire \myifu/myicache/_0586_ ;
wire \myifu/myicache/_0587_ ;
wire \myifu/myicache/_0588_ ;
wire \myifu/myicache/_0589_ ;
wire \myifu/myicache/_0590_ ;
wire \myifu/myicache/_0591_ ;
wire \myifu/myicache/_0592_ ;
wire \myifu/myicache/_0593_ ;
wire \myifu/myicache/_0594_ ;
wire \myifu/myicache/_0595_ ;
wire \myifu/myicache/_0596_ ;
wire \myifu/myicache/_0597_ ;
wire \myifu/myicache/_0598_ ;
wire \myifu/myicache/_0599_ ;
wire \myifu/myicache/_0600_ ;
wire \myifu/myicache/_0601_ ;
wire \myifu/myicache/_0602_ ;
wire \myifu/myicache/_0603_ ;
wire \myifu/myicache/_0604_ ;
wire \myifu/myicache/_0605_ ;
wire \myifu/myicache/_0606_ ;
wire \myifu/myicache/_0607_ ;
wire \myifu/myicache/_0608_ ;
wire \myifu/myicache/_0609_ ;
wire \myifu/myicache/_0610_ ;
wire \myifu/myicache/_0611_ ;
wire \myifu/myicache/_0612_ ;
wire \myifu/myicache/_0613_ ;
wire \myifu/myicache/_0614_ ;
wire \myifu/myicache/_0615_ ;
wire \myifu/myicache/_0616_ ;
wire \myifu/myicache/_0617_ ;
wire \myifu/myicache/_0618_ ;
wire \myifu/myicache/_0619_ ;
wire \myifu/myicache/_0620_ ;
wire \myifu/myicache/_0621_ ;
wire \myifu/myicache/_0622_ ;
wire \myifu/myicache/_0623_ ;
wire \myifu/myicache/_0624_ ;
wire \myifu/myicache/_0625_ ;
wire \myifu/myicache/_0626_ ;
wire \myifu/myicache/_0627_ ;
wire \myifu/myicache/_0628_ ;
wire \myifu/myicache/_0629_ ;
wire \myifu/myicache/_0630_ ;
wire \myifu/myicache/_0631_ ;
wire \myifu/myicache/_0632_ ;
wire \myifu/myicache/_0633_ ;
wire \myifu/myicache/_0634_ ;
wire \myifu/myicache/_0635_ ;
wire \myifu/myicache/_0636_ ;
wire \myifu/myicache/_0637_ ;
wire \myifu/myicache/_0638_ ;
wire \myifu/myicache/_0639_ ;
wire \myifu/myicache/_0640_ ;
wire \myifu/myicache/_0641_ ;
wire \myifu/myicache/_0642_ ;
wire \myifu/myicache/_0643_ ;
wire \myifu/myicache/_0644_ ;
wire \myifu/myicache/_0645_ ;
wire \myifu/myicache/_0646_ ;
wire \myifu/myicache/_0647_ ;
wire \myifu/myicache/_0648_ ;
wire \myifu/myicache/_0649_ ;
wire \myifu/myicache/_0650_ ;
wire \myifu/myicache/_0651_ ;
wire \myifu/myicache/_0652_ ;
wire \myifu/myicache/_0653_ ;
wire \myifu/myicache/_0654_ ;
wire \myifu/myicache/_0655_ ;
wire \myifu/myicache/_0656_ ;
wire \myifu/myicache/_0657_ ;
wire \myifu/myicache/_0658_ ;
wire \myifu/myicache/_0659_ ;
wire \myifu/myicache/_0660_ ;
wire \myifu/myicache/_0661_ ;
wire \myifu/myicache/_0662_ ;
wire \myifu/myicache/_0663_ ;
wire \myifu/myicache/_0664_ ;
wire \myifu/myicache/_0665_ ;
wire \myifu/myicache/_0666_ ;
wire \myifu/myicache/_0667_ ;
wire \myifu/myicache/_0668_ ;
wire \myifu/myicache/_0669_ ;
wire \myifu/myicache/_0670_ ;
wire \myifu/myicache/_0671_ ;
wire \myifu/myicache/_0672_ ;
wire \myifu/myicache/_0673_ ;
wire \myifu/myicache/_0674_ ;
wire \myifu/myicache/_0675_ ;
wire \myifu/myicache/_0676_ ;
wire \myifu/myicache/_0677_ ;
wire \myifu/myicache/_0678_ ;
wire \myifu/myicache/_0679_ ;
wire \myifu/myicache/_0680_ ;
wire \myifu/myicache/_0681_ ;
wire \myifu/myicache/_0682_ ;
wire \myifu/myicache/_0683_ ;
wire \myifu/myicache/_0684_ ;
wire \myifu/myicache/_0685_ ;
wire \myifu/myicache/_0686_ ;
wire \myifu/myicache/_0687_ ;
wire \myifu/myicache/_0688_ ;
wire \myifu/myicache/_0689_ ;
wire \myifu/myicache/_0690_ ;
wire \myifu/myicache/_0691_ ;
wire \myifu/myicache/_0692_ ;
wire \myifu/myicache/_0693_ ;
wire \myifu/myicache/_0694_ ;
wire \myifu/myicache/_0695_ ;
wire \myifu/myicache/_0696_ ;
wire \myifu/myicache/_0697_ ;
wire \myifu/myicache/_0698_ ;
wire \myifu/myicache/_0699_ ;
wire \myifu/myicache/_0700_ ;
wire \myifu/myicache/_0701_ ;
wire \myifu/myicache/_0702_ ;
wire \myifu/myicache/_0703_ ;
wire \myifu/myicache/_0704_ ;
wire \myifu/myicache/_0705_ ;
wire \myifu/myicache/_0706_ ;
wire \myifu/myicache/_0707_ ;
wire \myifu/myicache/_0708_ ;
wire \myifu/myicache/_0709_ ;
wire \myifu/myicache/_0710_ ;
wire \myifu/myicache/_0711_ ;
wire \myifu/myicache/_0712_ ;
wire \myifu/myicache/_0713_ ;
wire \myifu/myicache/_0714_ ;
wire \myifu/myicache/_0715_ ;
wire \myifu/myicache/_0716_ ;
wire \myifu/myicache/_0717_ ;
wire \myifu/myicache/_0718_ ;
wire \myifu/myicache/_0719_ ;
wire \myifu/myicache/_0720_ ;
wire \myifu/myicache/_0721_ ;
wire \myifu/myicache/_0722_ ;
wire \myifu/myicache/_0723_ ;
wire \myifu/myicache/_0724_ ;
wire \myifu/myicache/_0725_ ;
wire \myifu/myicache/_0726_ ;
wire \myifu/myicache/_0727_ ;
wire \myifu/myicache/_0728_ ;
wire \myifu/myicache/_0729_ ;
wire \myifu/myicache/_0730_ ;
wire \myifu/myicache/_0731_ ;
wire \myifu/myicache/_0732_ ;
wire \myifu/myicache/_0733_ ;
wire \myifu/myicache/_0734_ ;
wire \myifu/myicache/_0735_ ;
wire \myifu/myicache/_0736_ ;
wire \myifu/myicache/_0737_ ;
wire \myifu/myicache/_0738_ ;
wire \myifu/myicache/_0739_ ;
wire \myifu/myicache/_0740_ ;
wire \myifu/myicache/_0741_ ;
wire \myifu/myicache/_0742_ ;
wire \myifu/myicache/_0743_ ;
wire \myifu/myicache/_0744_ ;
wire \myifu/myicache/_0745_ ;
wire \myifu/myicache/_0746_ ;
wire \myifu/myicache/_0747_ ;
wire \myifu/myicache/_0748_ ;
wire \myifu/myicache/_0749_ ;
wire \myifu/myicache/_0750_ ;
wire \myifu/myicache/_0751_ ;
wire \myifu/myicache/_0752_ ;
wire \myifu/myicache/_0753_ ;
wire \myifu/myicache/_0754_ ;
wire \myifu/myicache/_0755_ ;
wire \myifu/myicache/_0756_ ;
wire \myifu/myicache/_0757_ ;
wire \myifu/myicache/_0758_ ;
wire \myifu/myicache/_0759_ ;
wire \myifu/myicache/_0760_ ;
wire \myifu/myicache/_0761_ ;
wire \myifu/myicache/_0762_ ;
wire \myifu/myicache/_0763_ ;
wire \myifu/myicache/_0764_ ;
wire \myifu/myicache/_0765_ ;
wire \myifu/myicache/_0766_ ;
wire \myifu/myicache/_0767_ ;
wire \myifu/myicache/_0768_ ;
wire \myifu/myicache/_0769_ ;
wire \myifu/myicache/_0770_ ;
wire \myifu/myicache/_0771_ ;
wire \myifu/myicache/_0772_ ;
wire \myifu/myicache/_0773_ ;
wire \myifu/myicache/_0774_ ;
wire \myifu/myicache/_0775_ ;
wire \myifu/myicache/_0776_ ;
wire \myifu/myicache/_0777_ ;
wire \myifu/myicache/_0778_ ;
wire \myifu/myicache/_0779_ ;
wire \myifu/myicache/_0780_ ;
wire \myifu/myicache/_0781_ ;
wire \myifu/myicache/_0782_ ;
wire \myifu/myicache/_0783_ ;
wire \myifu/myicache/_0784_ ;
wire \myifu/myicache/_0785_ ;
wire \myifu/myicache/_0786_ ;
wire \myifu/myicache/_0787_ ;
wire \myifu/myicache/_0788_ ;
wire \myifu/myicache/_0789_ ;
wire \myifu/myicache/_0790_ ;
wire \myifu/myicache/_0791_ ;
wire \myifu/myicache/_0792_ ;
wire \myifu/myicache/_0793_ ;
wire \myifu/myicache/_0794_ ;
wire \myifu/myicache/_0795_ ;
wire \myifu/myicache/_0796_ ;
wire \myifu/myicache/_0797_ ;
wire \myifu/myicache/_0798_ ;
wire \myifu/myicache/_0799_ ;
wire \myifu/myicache/_0800_ ;
wire \myifu/myicache/_0801_ ;
wire \myifu/myicache/_0802_ ;
wire \myifu/myicache/_0803_ ;
wire \myifu/myicache/_0804_ ;
wire \myifu/myicache/_0805_ ;
wire \myifu/myicache/_0806_ ;
wire \myifu/myicache/_0807_ ;
wire \myifu/myicache/_0808_ ;
wire \myifu/myicache/_0809_ ;
wire \myifu/myicache/_0810_ ;
wire \myifu/myicache/_0811_ ;
wire \myifu/myicache/_0812_ ;
wire \myifu/myicache/_0813_ ;
wire \myifu/myicache/_0814_ ;
wire \myifu/myicache/_0815_ ;
wire \myifu/myicache/_0816_ ;
wire \myifu/myicache/_0817_ ;
wire \myifu/myicache/_0818_ ;
wire \myifu/myicache/_0819_ ;
wire \myifu/myicache/_0820_ ;
wire \myifu/myicache/_0821_ ;
wire \myifu/myicache/_0822_ ;
wire \myifu/myicache/_0823_ ;
wire \myifu/myicache/_0824_ ;
wire \myifu/myicache/_0825_ ;
wire \myifu/myicache/_0826_ ;
wire \myifu/myicache/_0827_ ;
wire \myifu/myicache/_0828_ ;
wire \myifu/myicache/_0829_ ;
wire \myifu/myicache/_0830_ ;
wire \myifu/myicache/_0831_ ;
wire \myifu/myicache/_0832_ ;
wire \myifu/myicache/_0833_ ;
wire \myifu/myicache/_0834_ ;
wire \myifu/myicache/_0835_ ;
wire \myifu/myicache/_0836_ ;
wire \myifu/myicache/_0837_ ;
wire \myifu/myicache/_0838_ ;
wire \myifu/myicache/_0839_ ;
wire \myifu/myicache/_0840_ ;
wire \myifu/myicache/_0841_ ;
wire \myifu/myicache/_0842_ ;
wire \myifu/myicache/_0843_ ;
wire \myifu/myicache/_0844_ ;
wire \myifu/myicache/_0845_ ;
wire \myifu/myicache/_0846_ ;
wire \myifu/myicache/_0847_ ;
wire \myifu/myicache/_0848_ ;
wire \myifu/myicache/_0849_ ;
wire \myifu/myicache/_0850_ ;
wire \myifu/myicache/_0851_ ;
wire \myifu/myicache/_0852_ ;
wire \myifu/myicache/_0853_ ;
wire \myifu/myicache/_0854_ ;
wire \myifu/myicache/_0855_ ;
wire \myifu/myicache/_0856_ ;
wire \myifu/myicache/_0857_ ;
wire \myifu/myicache/_0858_ ;
wire \myifu/myicache/_0859_ ;
wire \myifu/myicache/_0860_ ;
wire \myifu/myicache/_0861_ ;
wire \myifu/myicache/_0862_ ;
wire \myifu/myicache/_0863_ ;
wire \myifu/myicache/_0864_ ;
wire \myifu/myicache/_0865_ ;
wire \myifu/myicache/_0866_ ;
wire \myifu/myicache/_0867_ ;
wire \myifu/myicache/_0868_ ;
wire \myifu/myicache/_0869_ ;
wire \myifu/myicache/_0870_ ;
wire \myifu/myicache/_0871_ ;
wire \myifu/myicache/_0872_ ;
wire \myifu/myicache/_0873_ ;
wire \myifu/myicache/_0874_ ;
wire \myifu/myicache/_0875_ ;
wire \myifu/myicache/_0876_ ;
wire \myifu/myicache/_0877_ ;
wire \myifu/myicache/_0878_ ;
wire \myifu/myicache/_0879_ ;
wire \myifu/myicache/_0880_ ;
wire \myifu/myicache/_0881_ ;
wire \myifu/myicache/_0882_ ;
wire \myifu/myicache/_0883_ ;
wire \myifu/myicache/_0884_ ;
wire \myifu/myicache/_0885_ ;
wire \myifu/myicache/_0886_ ;
wire \myifu/myicache/_0887_ ;
wire \myifu/myicache/_0888_ ;
wire \myifu/myicache/_0889_ ;
wire \myifu/myicache/_0890_ ;
wire \myifu/myicache/_0891_ ;
wire \myifu/myicache/_0892_ ;
wire \myifu/myicache/_0893_ ;
wire \myifu/myicache/_0894_ ;
wire \myifu/myicache/_0895_ ;
wire \myifu/myicache/_0896_ ;
wire \myifu/myicache/_0897_ ;
wire \myifu/myicache/_0898_ ;
wire \myifu/myicache/_0899_ ;
wire \myifu/myicache/_0900_ ;
wire \myifu/myicache/_0901_ ;
wire \myifu/myicache/_0902_ ;
wire \myifu/myicache/_0903_ ;
wire \myifu/myicache/_0904_ ;
wire \myifu/myicache/_0905_ ;
wire \myifu/myicache/_0906_ ;
wire \myifu/myicache/_0907_ ;
wire \myifu/myicache/_0908_ ;
wire \myifu/myicache/_0909_ ;
wire \myifu/myicache/_0910_ ;
wire \myifu/myicache/_0911_ ;
wire \myifu/myicache/_0912_ ;
wire \myifu/myicache/_0913_ ;
wire \myifu/myicache/_0914_ ;
wire \myifu/myicache/_0915_ ;
wire \myifu/myicache/_0916_ ;
wire \myifu/myicache/_0917_ ;
wire \myifu/myicache/_0918_ ;
wire \myifu/myicache/_0919_ ;
wire \myifu/myicache/_0920_ ;
wire \myifu/myicache/_0921_ ;
wire \myifu/myicache/_0922_ ;
wire \myifu/myicache/_0923_ ;
wire \myifu/myicache/_0924_ ;
wire \myifu/myicache/_0925_ ;
wire \myifu/myicache/_0926_ ;
wire \myifu/myicache/_0927_ ;
wire \myifu/myicache/_0928_ ;
wire \myifu/myicache/_0929_ ;
wire \myifu/myicache/_0930_ ;
wire \myifu/myicache/_0931_ ;
wire \myifu/myicache/_0932_ ;
wire \myifu/myicache/_0933_ ;
wire \myifu/myicache/_0934_ ;
wire \myifu/myicache/_0935_ ;
wire \myifu/myicache/_0936_ ;
wire \myifu/myicache/_0937_ ;
wire \myifu/myicache/_0938_ ;
wire \myifu/myicache/_0939_ ;
wire \myifu/myicache/_0940_ ;
wire \myifu/myicache/_0941_ ;
wire \myifu/myicache/_0942_ ;
wire \myifu/myicache/_0943_ ;
wire \myifu/myicache/_0944_ ;
wire \myifu/myicache/_0945_ ;
wire \myifu/myicache/_0946_ ;
wire \myifu/myicache/_0947_ ;
wire \myifu/myicache/_0948_ ;
wire \myifu/myicache/_0949_ ;
wire \myifu/myicache/_0950_ ;
wire \myifu/myicache/_0951_ ;
wire \myifu/myicache/_0952_ ;
wire \myifu/myicache/_0953_ ;
wire \myifu/myicache/_0954_ ;
wire \myifu/myicache/_0955_ ;
wire \myifu/myicache/_0956_ ;
wire \myifu/myicache/_0957_ ;
wire \myifu/myicache/_0958_ ;
wire \myifu/myicache/_0959_ ;
wire \myifu/myicache/_0960_ ;
wire \myifu/myicache/_0961_ ;
wire \myifu/myicache/_0962_ ;
wire \myifu/myicache/_0963_ ;
wire \myifu/myicache/_0964_ ;
wire \myifu/myicache/_0965_ ;
wire \myifu/myicache/_0966_ ;
wire \myifu/myicache/_0967_ ;
wire \myifu/myicache/_0968_ ;
wire \myifu/myicache/_0969_ ;
wire \myifu/myicache/_0970_ ;
wire \myifu/myicache/_0971_ ;
wire \myifu/myicache/_0972_ ;
wire \myifu/myicache/_0973_ ;
wire \myifu/myicache/_0974_ ;
wire \myifu/myicache/_0975_ ;
wire \myifu/myicache/_0976_ ;
wire \myifu/myicache/_0977_ ;
wire \myifu/myicache/_0978_ ;
wire \myifu/myicache/_0979_ ;
wire \myifu/myicache/_0980_ ;
wire \myifu/myicache/_0981_ ;
wire \myifu/myicache/_0982_ ;
wire \myifu/myicache/_0983_ ;
wire \myifu/myicache/_0984_ ;
wire \myifu/myicache/_0985_ ;
wire \myifu/myicache/_0986_ ;
wire \myifu/myicache/_0987_ ;
wire \myifu/myicache/_0988_ ;
wire \myifu/myicache/_0989_ ;
wire \myifu/myicache/_0990_ ;
wire \myifu/myicache/_0991_ ;
wire \myifu/myicache/_0992_ ;
wire \myifu/myicache/_0993_ ;
wire \myifu/myicache/_0994_ ;
wire \myifu/myicache/_0995_ ;
wire \myifu/myicache/_0996_ ;
wire \myifu/myicache/_0997_ ;
wire \myifu/myicache/_0998_ ;
wire \myifu/myicache/_0999_ ;
wire \myifu/myicache/_1000_ ;
wire \myifu/myicache/_1001_ ;
wire \myifu/myicache/_1002_ ;
wire \myifu/myicache/_1003_ ;
wire \myifu/myicache/_1004_ ;
wire \myifu/myicache/_1005_ ;
wire \myifu/myicache/_1006_ ;
wire \myifu/myicache/_1007_ ;
wire \myifu/myicache/_1008_ ;
wire \myifu/myicache/_1009_ ;
wire \myifu/myicache/_1010_ ;
wire \myifu/myicache/_1011_ ;
wire \myifu/myicache/_1012_ ;
wire \myifu/myicache/_1013_ ;
wire \myifu/myicache/_1014_ ;
wire \myifu/myicache/_1015_ ;
wire \myifu/myicache/_1016_ ;
wire \myifu/myicache/_1017_ ;
wire \myifu/myicache/_1018_ ;
wire \myifu/myicache/_1019_ ;
wire \myifu/myicache/_1020_ ;
wire \myifu/myicache/_1021_ ;
wire \myifu/myicache/_1022_ ;
wire \myifu/myicache/_1023_ ;
wire \myifu/myicache/_1024_ ;
wire \myifu/myicache/_1025_ ;
wire \myifu/myicache/_1026_ ;
wire \myifu/myicache/_1027_ ;
wire \myifu/myicache/_1028_ ;
wire \myifu/myicache/_1029_ ;
wire \myifu/myicache/_1030_ ;
wire \myifu/myicache/_1031_ ;
wire \myifu/myicache/_1032_ ;
wire \myifu/myicache/_1033_ ;
wire \myifu/myicache/_1034_ ;
wire \myifu/myicache/_1035_ ;
wire \myifu/myicache/_1036_ ;
wire \myifu/myicache/_1037_ ;
wire \myifu/myicache/_1038_ ;
wire \myifu/myicache/_1039_ ;
wire \myifu/myicache/_1040_ ;
wire \myifu/myicache/_1041_ ;
wire \myifu/myicache/_1042_ ;
wire \myifu/myicache/_1043_ ;
wire \myifu/myicache/_1044_ ;
wire \myifu/myicache/_1045_ ;
wire \myifu/myicache/_1046_ ;
wire \myifu/myicache/_1047_ ;
wire \myifu/myicache/_1048_ ;
wire \myifu/myicache/_1049_ ;
wire \myifu/myicache/_1050_ ;
wire \myifu/myicache/_1051_ ;
wire \myifu/myicache/_1052_ ;
wire \myifu/myicache/_1053_ ;
wire \myifu/myicache/_1054_ ;
wire \myifu/myicache/_1055_ ;
wire \myifu/myicache/_1056_ ;
wire \myifu/myicache/_1057_ ;
wire \myifu/myicache/_1058_ ;
wire \myifu/myicache/_1059_ ;
wire \myifu/myicache/_1060_ ;
wire \myifu/myicache/_1061_ ;
wire \myifu/myicache/_1062_ ;
wire \myifu/myicache/_1063_ ;
wire \myifu/myicache/_1064_ ;
wire \myifu/myicache/_1065_ ;
wire \myifu/myicache/_1066_ ;
wire \myifu/myicache/_1067_ ;
wire \myifu/myicache/_1068_ ;
wire \myifu/myicache/_1069_ ;
wire \myifu/myicache/_1070_ ;
wire \myifu/myicache/_1071_ ;
wire \myifu/myicache/_1072_ ;
wire \myifu/myicache/_1073_ ;
wire \myifu/myicache/_1074_ ;
wire \myifu/myicache/_1075_ ;
wire \myifu/myicache/_1076_ ;
wire \myifu/myicache/_1077_ ;
wire \myifu/myicache/_1078_ ;
wire \myifu/myicache/_1079_ ;
wire \myifu/myicache/_1080_ ;
wire \myifu/myicache/_1081_ ;
wire \myifu/myicache/_1082_ ;
wire \myifu/myicache/_1083_ ;
wire \myifu/myicache/_1084_ ;
wire \myifu/myicache/_1085_ ;
wire \myifu/myicache/_1086_ ;
wire \myifu/myicache/_1087_ ;
wire \myifu/myicache/_1088_ ;
wire \myifu/myicache/_1089_ ;
wire \myifu/myicache/_1090_ ;
wire \myifu/myicache/_1091_ ;
wire \myifu/myicache/_1092_ ;
wire \myifu/myicache/_1093_ ;
wire \myifu/myicache/_1094_ ;
wire \myifu/myicache/_1095_ ;
wire \myifu/myicache/_1096_ ;
wire \myifu/myicache/_1097_ ;
wire \myifu/myicache/_1098_ ;
wire \myifu/myicache/_1099_ ;
wire \myifu/myicache/_1100_ ;
wire \myifu/myicache/_1101_ ;
wire \myifu/myicache/_1102_ ;
wire \myifu/myicache/_1103_ ;
wire \myifu/myicache/_1104_ ;
wire \myifu/myicache/_1105_ ;
wire \myifu/myicache/_1106_ ;
wire \myifu/myicache/_1107_ ;
wire \myifu/myicache/_1108_ ;
wire \myifu/myicache/_1109_ ;
wire \myifu/myicache/_1110_ ;
wire \myifu/myicache/_1111_ ;
wire \myifu/myicache/_1112_ ;
wire \myifu/myicache/_1113_ ;
wire \myifu/myicache/_1114_ ;
wire \myifu/myicache/_1115_ ;
wire \myifu/myicache/_1116_ ;
wire \myifu/myicache/_1117_ ;
wire \myifu/myicache/_1118_ ;
wire \myifu/myicache/_1119_ ;
wire \myifu/myicache/_1120_ ;
wire \myifu/myicache/_1121_ ;
wire \myifu/myicache/_1122_ ;
wire \myifu/myicache/_1123_ ;
wire \myifu/myicache/_1124_ ;
wire \myifu/myicache/_1125_ ;
wire \myifu/myicache/_1126_ ;
wire \myifu/myicache/_1127_ ;
wire \myifu/myicache/_1128_ ;
wire \myifu/myicache/_1129_ ;
wire \myifu/myicache/_1130_ ;
wire \myifu/myicache/_1131_ ;
wire \myifu/myicache/_1132_ ;
wire \myifu/myicache/_1133_ ;
wire \myifu/myicache/_1134_ ;
wire \myifu/myicache/_1135_ ;
wire \myifu/myicache/_1136_ ;
wire \myifu/myicache/_1137_ ;
wire \myifu/myicache/_1138_ ;
wire \myifu/myicache/_1139_ ;
wire \myifu/myicache/_1140_ ;
wire \myifu/myicache/_1141_ ;
wire \myifu/myicache/_1142_ ;
wire \myifu/myicache/_1143_ ;
wire \myifu/myicache/_1144_ ;
wire \myifu/myicache/_1145_ ;
wire \myifu/myicache/_1146_ ;
wire \myifu/myicache/_1147_ ;
wire \myifu/myicache/_1148_ ;
wire \myifu/myicache/_1149_ ;
wire \myifu/myicache/_1150_ ;
wire \myifu/myicache/_1151_ ;
wire \myifu/myicache/_1152_ ;
wire \myifu/myicache/_1153_ ;
wire \myifu/myicache/_1154_ ;
wire \myifu/myicache/_1155_ ;
wire \myifu/myicache/_1156_ ;
wire \myifu/myicache/_1157_ ;
wire \myifu/myicache/_1158_ ;
wire \myifu/myicache/_1159_ ;
wire \myifu/myicache/_1160_ ;
wire \myifu/myicache/_1161_ ;
wire \myifu/myicache/_1162_ ;
wire \myifu/myicache/_1163_ ;
wire \myifu/myicache/_1164_ ;
wire \myifu/myicache/_1165_ ;
wire \myifu/myicache/_1166_ ;
wire \myifu/myicache/_1167_ ;
wire \myifu/myicache/_1168_ ;
wire \myifu/myicache/_1169_ ;
wire \myifu/myicache/_1170_ ;
wire \myifu/myicache/_1171_ ;
wire \myifu/myicache/_1172_ ;
wire \myifu/myicache/_1173_ ;
wire \myifu/myicache/_1174_ ;
wire \myifu/myicache/_1175_ ;
wire \myifu/myicache/_1176_ ;
wire \myifu/myicache/_1177_ ;
wire \myifu/myicache/_1178_ ;
wire \myifu/myicache/_1179_ ;
wire \myifu/myicache/_1180_ ;
wire \myifu/myicache/_1181_ ;
wire \myifu/myicache/_1182_ ;
wire \myifu/myicache/_1183_ ;
wire \myifu/myicache/_1184_ ;
wire \myifu/myicache/_1185_ ;
wire \myifu/myicache/_1186_ ;
wire \myifu/myicache/_1187_ ;
wire \myifu/myicache/_1188_ ;
wire \myifu/myicache/_1189_ ;
wire \myifu/myicache/_1190_ ;
wire \myifu/myicache/_1191_ ;
wire \myifu/myicache/_1192_ ;
wire \myifu/myicache/_1193_ ;
wire \myifu/myicache/_1194_ ;
wire \myifu/myicache/_1195_ ;
wire \myifu/myicache/_1196_ ;
wire \myifu/myicache/_1197_ ;
wire \myifu/myicache/_1198_ ;
wire \myifu/myicache/_1199_ ;
wire \myifu/myicache/_1200_ ;
wire \myifu/myicache/_1201_ ;
wire \myifu/myicache/_1202_ ;
wire \myifu/myicache/_1203_ ;
wire \myifu/myicache/_1204_ ;
wire \myifu/myicache/_1205_ ;
wire \myifu/myicache/_1206_ ;
wire \myifu/myicache/_1207_ ;
wire \myifu/myicache/_1208_ ;
wire \myifu/myicache/_1209_ ;
wire \myifu/myicache/_1210_ ;
wire \myifu/myicache/_1211_ ;
wire \myifu/myicache/_1212_ ;
wire \myifu/myicache/_1213_ ;
wire \myifu/myicache/_1214_ ;
wire \myifu/myicache/_1215_ ;
wire \myifu/myicache/_1216_ ;
wire \myifu/myicache/_1217_ ;
wire \myifu/myicache/_1218_ ;
wire \myifu/myicache/_1219_ ;
wire \myifu/myicache/_1220_ ;
wire \myifu/myicache/_1221_ ;
wire \myifu/myicache/_1222_ ;
wire \myifu/myicache/_1223_ ;
wire \myifu/myicache/_1224_ ;
wire \myifu/myicache/_1225_ ;
wire \myifu/myicache/_1226_ ;
wire \myifu/myicache/_1227_ ;
wire \myifu/myicache/_1228_ ;
wire \myifu/myicache/_1229_ ;
wire \myifu/myicache/_1230_ ;
wire \myifu/myicache/_1231_ ;
wire \myifu/myicache/_1232_ ;
wire \myifu/myicache/_1233_ ;
wire \myifu/myicache/_1234_ ;
wire \myifu/myicache/_1235_ ;
wire \myifu/myicache/_1236_ ;
wire \myifu/myicache/_1237_ ;
wire \myifu/myicache/_1238_ ;
wire \myifu/myicache/_1239_ ;
wire \myifu/myicache/_1240_ ;
wire \myifu/myicache/_1241_ ;
wire \myifu/myicache/_1242_ ;
wire \myifu/myicache/_1243_ ;
wire \myifu/myicache/_1244_ ;
wire \myifu/myicache/_1245_ ;
wire \myifu/myicache/_1246_ ;
wire \myifu/myicache/_1247_ ;
wire \myifu/myicache/_1248_ ;
wire \myifu/myicache/_1249_ ;
wire \myifu/myicache/_1250_ ;
wire \myifu/myicache/_1251_ ;
wire \myifu/myicache/_1252_ ;
wire \myifu/myicache/_1253_ ;
wire \myifu/myicache/_1254_ ;
wire \myifu/myicache/_1255_ ;
wire \myifu/myicache/_1256_ ;
wire \myifu/myicache/_1257_ ;
wire \myifu/myicache/_1258_ ;
wire \myifu/myicache/_1259_ ;
wire \myifu/myicache/_1260_ ;
wire \myifu/myicache/_1261_ ;
wire \myifu/myicache/_1262_ ;
wire \myifu/myicache/_1263_ ;
wire \myifu/myicache/_1264_ ;
wire \myifu/myicache/_1265_ ;
wire \myifu/myicache/_1266_ ;
wire \myifu/myicache/_1267_ ;
wire \myifu/myicache/_1268_ ;
wire \myifu/myicache/_1269_ ;
wire \myifu/myicache/_1270_ ;
wire \myifu/myicache/_1271_ ;
wire \myifu/myicache/_1272_ ;
wire \myifu/myicache/_1273_ ;
wire \myifu/myicache/_1274_ ;
wire \myifu/myicache/_1275_ ;
wire \myifu/myicache/_1276_ ;
wire \myifu/myicache/_1277_ ;
wire \myifu/myicache/_1278_ ;
wire \myifu/myicache/_1279_ ;
wire \myifu/myicache/_1280_ ;
wire \myifu/myicache/_1281_ ;
wire \myifu/myicache/_1282_ ;
wire \myifu/myicache/_1283_ ;
wire \myifu/myicache/_1284_ ;
wire \myifu/myicache/_1285_ ;
wire \myifu/myicache/_1286_ ;
wire \myifu/myicache/_1287_ ;
wire \myifu/myicache/_1288_ ;
wire \myifu/myicache/_1289_ ;
wire \myifu/myicache/_1290_ ;
wire \myifu/myicache/_1291_ ;
wire \myifu/myicache/_1292_ ;
wire \myifu/myicache/_1293_ ;
wire \myifu/myicache/_1294_ ;
wire \myifu/myicache/_1295_ ;
wire \myifu/myicache/_1296_ ;
wire \myifu/myicache/_1297_ ;
wire \myifu/myicache/_1298_ ;
wire \myifu/myicache/_1299_ ;
wire \myifu/myicache/_1300_ ;
wire \myifu/myicache/_1301_ ;
wire \myifu/myicache/_1302_ ;
wire \myifu/myicache/_1303_ ;
wire \myifu/myicache/_1304_ ;
wire \myifu/myicache/_1305_ ;
wire \myifu/myicache/_1306_ ;
wire \myifu/myicache/_1307_ ;
wire \myifu/myicache/_1308_ ;
wire \myifu/myicache/_1309_ ;
wire \myifu/myicache/_1310_ ;
wire \myifu/myicache/_1311_ ;
wire \myifu/myicache/_1312_ ;
wire \myifu/myicache/_1313_ ;
wire \myifu/myicache/_1314_ ;
wire \myifu/myicache/_1315_ ;
wire \myifu/myicache/_1316_ ;
wire \myifu/myicache/_1317_ ;
wire \myifu/myicache/_1318_ ;
wire \myifu/myicache/_1319_ ;
wire \myifu/myicache/_1320_ ;
wire \myifu/myicache/_1321_ ;
wire \myifu/myicache/_1322_ ;
wire \myifu/myicache/_1323_ ;
wire \myifu/myicache/_1324_ ;
wire \myifu/myicache/_1325_ ;
wire \myifu/myicache/_1326_ ;
wire \myifu/myicache/_1327_ ;
wire \myifu/myicache/_1328_ ;
wire \myifu/myicache/_1329_ ;
wire \myifu/myicache/_1330_ ;
wire \myifu/myicache/_1331_ ;
wire \myifu/myicache/_1332_ ;
wire \myifu/myicache/_1333_ ;
wire \myifu/myicache/_1334_ ;
wire \myifu/myicache/_1335_ ;
wire \myifu/myicache/_1336_ ;
wire \myifu/myicache/_1337_ ;
wire \myifu/myicache/_1338_ ;
wire \myifu/myicache/_1339_ ;
wire \myifu/myicache/_1340_ ;
wire \myifu/myicache/_1341_ ;
wire \myifu/myicache/_1342_ ;
wire \myifu/myicache/_1343_ ;
wire \myifu/myicache/_1344_ ;
wire \myifu/myicache/_1345_ ;
wire \myifu/myicache/_1346_ ;
wire \myifu/myicache/_1347_ ;
wire \myifu/myicache/_1348_ ;
wire \myifu/myicache/_1349_ ;
wire \myifu/myicache/_1350_ ;
wire \myifu/myicache/_1351_ ;
wire \myifu/myicache/_1352_ ;
wire \myifu/myicache/_1353_ ;
wire \myifu/myicache/_1354_ ;
wire \myifu/myicache/_1355_ ;
wire \myifu/myicache/_1356_ ;
wire \myifu/myicache/_1357_ ;
wire \myifu/myicache/_1358_ ;
wire \myifu/myicache/_1359_ ;
wire \myifu/myicache/_1360_ ;
wire \myifu/myicache/_1361_ ;
wire \myifu/myicache/_1362_ ;
wire \myifu/myicache/_1363_ ;
wire \myifu/myicache/_1364_ ;
wire \myifu/myicache/_1365_ ;
wire \myifu/myicache/_1366_ ;
wire \myifu/myicache/_1367_ ;
wire \myifu/myicache/_1368_ ;
wire \myifu/myicache/_1369_ ;
wire \myifu/myicache/_1370_ ;
wire \myifu/myicache/_1371_ ;
wire \myifu/myicache/_1372_ ;
wire \myifu/myicache/_1373_ ;
wire \myifu/myicache/_1374_ ;
wire \myifu/myicache/_1375_ ;
wire \myifu/myicache/_1376_ ;
wire \myifu/myicache/_1377_ ;
wire \myifu/myicache/_1378_ ;
wire \myifu/myicache/_1379_ ;
wire \myifu/myicache/_1380_ ;
wire \myifu/myicache/_1381_ ;
wire \myifu/myicache/_1382_ ;
wire \myifu/myicache/_1383_ ;
wire \myifu/myicache/_1384_ ;
wire \myifu/myicache/_1385_ ;
wire \myifu/myicache/_1386_ ;
wire \myifu/myicache/_1387_ ;
wire \myifu/myicache/_1388_ ;
wire \myifu/myicache/_1389_ ;
wire \myifu/myicache/_1390_ ;
wire \myifu/myicache/_1391_ ;
wire \myifu/myicache/_1392_ ;
wire \myifu/myicache/_1393_ ;
wire \myifu/myicache/_1394_ ;
wire \myifu/myicache/_1395_ ;
wire \myifu/myicache/_1396_ ;
wire \myifu/myicache/_1397_ ;
wire \myifu/myicache/_1398_ ;
wire \myifu/myicache/_1399_ ;
wire \myifu/myicache/_1400_ ;
wire \myifu/myicache/_1401_ ;
wire \myifu/myicache/_1402_ ;
wire \myifu/myicache/_1403_ ;
wire \myifu/myicache/_1404_ ;
wire \myifu/myicache/_1405_ ;
wire \myifu/myicache/_1406_ ;
wire \myifu/myicache/_1407_ ;
wire \myifu/myicache/_1408_ ;
wire \myifu/myicache/_1409_ ;
wire \myifu/myicache/_1410_ ;
wire \myifu/myicache/_1411_ ;
wire \myifu/myicache/_1412_ ;
wire \myifu/myicache/_1413_ ;
wire \myifu/myicache/_1414_ ;
wire \myifu/myicache/_1415_ ;
wire \myifu/myicache/_1416_ ;
wire \myifu/myicache/_1417_ ;
wire \myifu/myicache/_1418_ ;
wire \myifu/myicache/_1419_ ;
wire \myifu/myicache/_1420_ ;
wire \myifu/myicache/_1421_ ;
wire \myifu/myicache/_1422_ ;
wire \myifu/myicache/_1423_ ;
wire \myifu/myicache/_1424_ ;
wire \myifu/myicache/_1425_ ;
wire \myifu/myicache/_1426_ ;
wire \myifu/myicache/_1427_ ;
wire \myifu/myicache/_1428_ ;
wire \myifu/myicache/_1429_ ;
wire \myifu/myicache/_1430_ ;
wire \myifu/myicache/_1431_ ;
wire \myifu/myicache/_1432_ ;
wire \myifu/myicache/_1433_ ;
wire \myifu/myicache/_1434_ ;
wire \myifu/myicache/_1435_ ;
wire \myifu/myicache/_1436_ ;
wire \myifu/myicache/_1437_ ;
wire \myifu/myicache/_1438_ ;
wire \myifu/myicache/_1439_ ;
wire \myifu/myicache/_1440_ ;
wire \myifu/myicache/_1441_ ;
wire \myifu/myicache/_1442_ ;
wire \myifu/myicache/_1443_ ;
wire \myifu/myicache/_1444_ ;
wire \myifu/myicache/_1445_ ;
wire \myifu/myicache/_1446_ ;
wire \myifu/myicache/_1447_ ;
wire \myifu/myicache/_1448_ ;
wire \myifu/myicache/_1449_ ;
wire \myifu/myicache/_1450_ ;
wire \myifu/myicache/_1451_ ;
wire \myifu/myicache/_1452_ ;
wire \myifu/myicache/_1453_ ;
wire \myifu/myicache/_1454_ ;
wire \myifu/myicache/_1455_ ;
wire \myifu/myicache/_1456_ ;
wire \myifu/myicache/_1457_ ;
wire \myifu/myicache/_1458_ ;
wire \myifu/myicache/_1459_ ;
wire \myifu/myicache/_1460_ ;
wire \myifu/myicache/_1461_ ;
wire \myifu/myicache/_1462_ ;
wire \myifu/myicache/_1463_ ;
wire \myifu/myicache/_1464_ ;
wire \myifu/myicache/_1465_ ;
wire \myifu/myicache/_1466_ ;
wire \myifu/myicache/_1467_ ;
wire \myifu/myicache/_1468_ ;
wire \myifu/myicache/_1469_ ;
wire \myifu/myicache/_1470_ ;
wire \myifu/myicache/_1471_ ;
wire \myifu/myicache/_1472_ ;
wire \myifu/myicache/_1473_ ;
wire \myifu/myicache/_1474_ ;
wire \myifu/myicache/_1475_ ;
wire \myifu/myicache/_1476_ ;
wire \myifu/myicache/_1477_ ;
wire \myifu/myicache/_1478_ ;
wire \myifu/myicache/_1479_ ;
wire \myifu/myicache/_1480_ ;
wire \myifu/myicache/_1481_ ;
wire \myifu/myicache/_1482_ ;
wire \myifu/myicache/_1483_ ;
wire \myifu/myicache/_1484_ ;
wire \myifu/myicache/_1485_ ;
wire \myifu/myicache/_1486_ ;
wire \myifu/myicache/_1487_ ;
wire \myifu/myicache/_1488_ ;
wire \myifu/myicache/_1489_ ;
wire \myifu/myicache/_1490_ ;
wire \myifu/myicache/_1491_ ;
wire \myifu/myicache/_1492_ ;
wire \myifu/myicache/_1493_ ;
wire \myifu/myicache/_1494_ ;
wire \myifu/myicache/_1495_ ;
wire \myifu/myicache/_1496_ ;
wire \myifu/myicache/_1497_ ;
wire \myifu/myicache/_1498_ ;
wire \myifu/myicache/_1499_ ;
wire \myifu/myicache/_1500_ ;
wire \myifu/myicache/_1501_ ;
wire \myifu/myicache/_1502_ ;
wire \myifu/myicache/_1503_ ;
wire \myifu/myicache/_1504_ ;
wire \myifu/myicache/_1505_ ;
wire \myifu/myicache/_1506_ ;
wire \myifu/myicache/_1507_ ;
wire \myifu/myicache/_1508_ ;
wire \myifu/myicache/_1509_ ;
wire \myifu/myicache/_1510_ ;
wire \myifu/myicache/_1511_ ;
wire \myifu/myicache/_1512_ ;
wire \myifu/myicache/_1513_ ;
wire \myifu/myicache/_1514_ ;
wire \myifu/myicache/_1515_ ;
wire \myifu/myicache/_1516_ ;
wire \myifu/myicache/_1517_ ;
wire \myifu/myicache/_1518_ ;
wire \myifu/myicache/_1519_ ;
wire \myifu/myicache/_1520_ ;
wire \myifu/myicache/_1521_ ;
wire \myifu/myicache/_1522_ ;
wire \myifu/myicache/_1523_ ;
wire \myifu/myicache/_1524_ ;
wire \myifu/myicache/_1525_ ;
wire \myifu/myicache/_1526_ ;
wire \myifu/myicache/_1527_ ;
wire \myifu/myicache/_1528_ ;
wire \myifu/myicache/_1529_ ;
wire \myifu/myicache/_1530_ ;
wire \myifu/myicache/_1531_ ;
wire \myifu/myicache/_1532_ ;
wire \myifu/myicache/_1533_ ;
wire \myifu/myicache/_1534_ ;
wire \myifu/myicache/_1535_ ;
wire \myifu/myicache/_1536_ ;
wire \myifu/myicache/_1537_ ;
wire \myifu/myicache/_1538_ ;
wire \myifu/myicache/_1539_ ;
wire \myifu/myicache/_1540_ ;
wire \myifu/myicache/_1541_ ;
wire \myifu/myicache/_1542_ ;
wire \myifu/myicache/_1543_ ;
wire \myifu/myicache/_1544_ ;
wire \myifu/myicache/_1545_ ;
wire \myifu/myicache/_1546_ ;
wire \myifu/myicache/_1547_ ;
wire \myifu/myicache/_1548_ ;
wire \myifu/myicache/_1549_ ;
wire \myifu/myicache/_1550_ ;
wire \myifu/myicache/_1551_ ;
wire \myifu/myicache/_1552_ ;
wire \myifu/myicache/_1553_ ;
wire \myifu/myicache/_1554_ ;
wire \myifu/myicache/_1555_ ;
wire \myifu/myicache/_1556_ ;
wire \myifu/myicache/_1557_ ;
wire \myifu/myicache/_1558_ ;
wire \myifu/myicache/_1559_ ;
wire \myifu/myicache/_1560_ ;
wire \myifu/myicache/_1561_ ;
wire \myifu/myicache/_1562_ ;
wire \myifu/myicache/_1563_ ;
wire \myifu/myicache/_1564_ ;
wire \myifu/myicache/_1565_ ;
wire \myifu/myicache/_1566_ ;
wire \myifu/myicache/_1567_ ;
wire \myifu/myicache/_1568_ ;
wire \myifu/myicache/_1569_ ;
wire \myifu/myicache/_1570_ ;
wire \myifu/myicache/_1571_ ;
wire \myifu/myicache/_1572_ ;
wire \myifu/myicache/_1573_ ;
wire \myifu/myicache/_1574_ ;
wire \myifu/myicache/_1575_ ;
wire \myifu/myicache/_1576_ ;
wire \myifu/myicache/_1577_ ;
wire \myifu/myicache/_1578_ ;
wire \myifu/myicache/_1579_ ;
wire \myifu/myicache/_1580_ ;
wire \myifu/myicache/_1581_ ;
wire \myifu/myicache/_1582_ ;
wire \myifu/myicache/_1583_ ;
wire \myifu/myicache/_1584_ ;
wire \myifu/myicache/_1585_ ;
wire \myifu/myicache/_1586_ ;
wire \myifu/myicache/_1587_ ;
wire \myifu/myicache/_1588_ ;
wire \myifu/myicache/_1589_ ;
wire \myifu/myicache/_1590_ ;
wire \myifu/myicache/_1591_ ;
wire \myifu/myicache/_1592_ ;
wire \myifu/myicache/_1593_ ;
wire \myifu/myicache/_1594_ ;
wire \myifu/myicache/_1595_ ;
wire \myifu/myicache/_1596_ ;
wire \myifu/myicache/_1597_ ;
wire \myifu/myicache/_1598_ ;
wire \myifu/myicache/_1599_ ;
wire \myifu/myicache/_1600_ ;
wire \myifu/myicache/_1601_ ;
wire \myifu/myicache/_1602_ ;
wire \myifu/myicache/_1603_ ;
wire \myifu/myicache/_1604_ ;
wire \myifu/myicache/_1605_ ;
wire \myifu/myicache/_1606_ ;
wire \myifu/myicache/_1607_ ;
wire \myifu/myicache/_1608_ ;
wire \myifu/myicache/_1609_ ;
wire \myifu/myicache/_1610_ ;
wire \myifu/myicache/_1611_ ;
wire \myifu/myicache/_1612_ ;
wire \myifu/myicache/_1613_ ;
wire \myifu/myicache/_1614_ ;
wire \myifu/myicache/_1615_ ;
wire \myifu/myicache/_1616_ ;
wire \myifu/myicache/_1617_ ;
wire \myifu/myicache/_1618_ ;
wire \myifu/myicache/_1619_ ;
wire \myifu/myicache/_1620_ ;
wire \myifu/myicache/_1621_ ;
wire \myifu/myicache/_1622_ ;
wire \myifu/myicache/_1623_ ;
wire \myifu/myicache/_1624_ ;
wire \myifu/myicache/_1625_ ;
wire \myifu/myicache/_1626_ ;
wire \myifu/myicache/_1627_ ;
wire \myifu/myicache/_1628_ ;
wire \myifu/myicache/_1629_ ;
wire \myifu/myicache/_1630_ ;
wire \myifu/myicache/_1631_ ;
wire \myifu/myicache/_1632_ ;
wire \myifu/myicache/_1633_ ;
wire \myifu/myicache/_1634_ ;
wire \myifu/myicache/_1635_ ;
wire \myifu/myicache/_1636_ ;
wire \myifu/myicache/_1637_ ;
wire \myifu/myicache/_1638_ ;
wire \myifu/myicache/_1639_ ;
wire \myifu/myicache/_1640_ ;
wire \myifu/myicache/_1641_ ;
wire \myifu/myicache/_1642_ ;
wire \myifu/myicache/_1643_ ;
wire \myifu/myicache/_1644_ ;
wire \myifu/myicache/_1645_ ;
wire \myifu/myicache/_1646_ ;
wire \myifu/myicache/_1647_ ;
wire \myifu/myicache/_1648_ ;
wire \myifu/myicache/_1649_ ;
wire \myifu/myicache/_1650_ ;
wire \myifu/myicache/_1651_ ;
wire \myifu/myicache/_1652_ ;
wire \myifu/myicache/_1653_ ;
wire \myifu/myicache/_1654_ ;
wire \myifu/myicache/_1655_ ;
wire \myifu/myicache/_1656_ ;
wire \myifu/myicache/_1657_ ;
wire \myifu/myicache/_1658_ ;
wire \myifu/myicache/_1659_ ;
wire \myifu/myicache/_1660_ ;
wire \myifu/myicache/_1661_ ;
wire \myifu/myicache/_1662_ ;
wire \myifu/myicache/_1663_ ;
wire \myifu/myicache/_1664_ ;
wire \myifu/myicache/_1665_ ;
wire \myifu/myicache/_1666_ ;
wire \myifu/myicache/_1667_ ;
wire \myifu/myicache/_1668_ ;
wire \myifu/myicache/_1669_ ;
wire \myifu/myicache/_1670_ ;
wire \myifu/myicache/_1671_ ;
wire \myifu/myicache/_1672_ ;
wire \myifu/myicache/_1673_ ;
wire \myifu/myicache/_1674_ ;
wire \myifu/myicache/_1675_ ;
wire \myifu/myicache/_1676_ ;
wire \myifu/myicache/_1677_ ;
wire \myifu/myicache/_1678_ ;
wire \myifu/myicache/_1679_ ;
wire \myifu/myicache/_1680_ ;
wire \myifu/myicache/_1681_ ;
wire \myifu/myicache/_1682_ ;
wire \myifu/myicache/_1683_ ;
wire \myifu/myicache/_1684_ ;
wire \myifu/myicache/_1685_ ;
wire \myifu/myicache/_1686_ ;
wire \myifu/myicache/_1687_ ;
wire \myifu/myicache/_1688_ ;
wire \myifu/myicache/_1689_ ;
wire \myifu/myicache/_1690_ ;
wire \myifu/myicache/_1691_ ;
wire \myifu/myicache/_1692_ ;
wire \myifu/myicache/_1693_ ;
wire \myifu/myicache/_1694_ ;
wire \myifu/myicache/_1695_ ;
wire \myifu/myicache/_1696_ ;
wire \myifu/myicache/_1697_ ;
wire \myifu/myicache/_1698_ ;
wire \myifu/myicache/_1699_ ;
wire \myifu/myicache/_1700_ ;
wire \myifu/myicache/_1701_ ;
wire \myifu/myicache/_1702_ ;
wire \myifu/myicache/_1703_ ;
wire \myifu/myicache/_1704_ ;
wire \myifu/myicache/_1705_ ;
wire \myifu/myicache/_1706_ ;
wire \myifu/myicache/_1707_ ;
wire \myifu/myicache/_1708_ ;
wire \myifu/myicache/_1709_ ;
wire \myifu/myicache/_1710_ ;
wire \myifu/myicache/_1711_ ;
wire \myifu/myicache/_1712_ ;
wire \myifu/myicache/_1713_ ;
wire \myifu/myicache/_1714_ ;
wire \myifu/myicache/_1715_ ;
wire \myifu/myicache/_1716_ ;
wire \myifu/myicache/_1717_ ;
wire \myifu/myicache/_1718_ ;
wire \myifu/myicache/_1719_ ;
wire \myifu/myicache/_1720_ ;
wire \myifu/myicache/_1721_ ;
wire \myifu/myicache/_1722_ ;
wire \myifu/myicache/_1723_ ;
wire \myifu/myicache/_1724_ ;
wire \myifu/myicache/_1725_ ;
wire \myifu/myicache/_1726_ ;
wire \myifu/myicache/_1727_ ;
wire \myifu/myicache/_1728_ ;
wire \myifu/myicache/_1729_ ;
wire \myifu/myicache/_1730_ ;
wire \myifu/myicache/_1731_ ;
wire \myifu/myicache/_1732_ ;
wire \myifu/myicache/_1733_ ;
wire \myifu/myicache/_1734_ ;
wire \myifu/myicache/_1735_ ;
wire \myifu/myicache/_1736_ ;
wire \myifu/myicache/_1737_ ;
wire \myifu/myicache/_1738_ ;
wire \myifu/myicache/_1739_ ;
wire \myifu/myicache/_1740_ ;
wire \myifu/myicache/_1741_ ;
wire \myifu/myicache/_1742_ ;
wire \myifu/myicache/_1743_ ;
wire \myifu/myicache/_1744_ ;
wire \myifu/myicache/_1745_ ;
wire \myifu/myicache/_1746_ ;
wire \myifu/myicache/_1747_ ;
wire \myifu/myicache/_1748_ ;
wire \myifu/myicache/_1749_ ;
wire \myifu/myicache/_1750_ ;
wire \myifu/myicache/_1751_ ;
wire \myifu/myicache/_1752_ ;
wire \myifu/myicache/_1753_ ;
wire \myifu/myicache/_1754_ ;
wire \myifu/myicache/_1755_ ;
wire \myifu/myicache/_1756_ ;
wire \myifu/myicache/_1757_ ;
wire \myifu/myicache/_1758_ ;
wire \myifu/myicache/_1759_ ;
wire \myifu/myicache/_1760_ ;
wire \myifu/myicache/_1761_ ;
wire \myifu/myicache/_1762_ ;
wire \myifu/myicache/_1763_ ;
wire \myifu/myicache/_1764_ ;
wire \myifu/myicache/_1765_ ;
wire \myifu/myicache/_1766_ ;
wire \myifu/myicache/_1767_ ;
wire \myifu/myicache/_1768_ ;
wire \myifu/myicache/_1769_ ;
wire \myifu/myicache/_1770_ ;
wire \myifu/myicache/_1771_ ;
wire \myifu/myicache/_1772_ ;
wire \myifu/myicache/_1773_ ;
wire \myifu/myicache/_1774_ ;
wire \myifu/myicache/_1775_ ;
wire \myifu/myicache/_1776_ ;
wire \myifu/myicache/_1777_ ;
wire \myifu/myicache/_1778_ ;
wire \myifu/myicache/_1779_ ;
wire \myifu/myicache/_1780_ ;
wire \myifu/myicache/_1781_ ;
wire \myifu/myicache/_1782_ ;
wire \myifu/myicache/_1783_ ;
wire \myifu/myicache/_1784_ ;
wire \myifu/myicache/_1785_ ;
wire \myifu/myicache/_1786_ ;
wire \myifu/myicache/_1787_ ;
wire \myifu/myicache/_1788_ ;
wire \myifu/myicache/_1789_ ;
wire \myifu/myicache/_1790_ ;
wire \myifu/myicache/_1791_ ;
wire \myifu/myicache/_1792_ ;
wire \myifu/myicache/_1793_ ;
wire \myifu/myicache/_1794_ ;
wire \myifu/myicache/_1795_ ;
wire \myifu/myicache/_1796_ ;
wire \myifu/myicache/_1797_ ;
wire \myifu/myicache/_1798_ ;
wire \myifu/myicache/_1799_ ;
wire \myifu/myicache/_1800_ ;
wire \myifu/myicache/_1801_ ;
wire \myifu/myicache/_1802_ ;
wire \myifu/myicache/_1803_ ;
wire \myifu/myicache/_1804_ ;
wire \myifu/myicache/_1805_ ;
wire \myifu/myicache/_1806_ ;
wire \myifu/myicache/_1807_ ;
wire \myifu/myicache/_1808_ ;
wire \myifu/myicache/_1809_ ;
wire \myifu/myicache/_1810_ ;
wire \myifu/myicache/_1811_ ;
wire \myifu/myicache/_1812_ ;
wire \myifu/myicache/_1813_ ;
wire \myifu/myicache/_1814_ ;
wire \myifu/myicache/_1815_ ;
wire \myifu/myicache/_1816_ ;
wire \myifu/myicache/_1817_ ;
wire \myifu/myicache/_1818_ ;
wire \myifu/myicache/_1819_ ;
wire \myifu/myicache/_1820_ ;
wire \myifu/myicache/_1821_ ;
wire \myifu/myicache/_1822_ ;
wire \myifu/myicache/_1823_ ;
wire \myifu/myicache/_1824_ ;
wire \myifu/myicache/_1825_ ;
wire \myifu/myicache/_1826_ ;
wire \myifu/myicache/_1827_ ;
wire \myifu/myicache/_1828_ ;
wire \myifu/myicache/_1829_ ;
wire \myifu/myicache/_1830_ ;
wire \myifu/myicache/_1831_ ;
wire \myifu/myicache/_1832_ ;
wire \myifu/myicache/_1833_ ;
wire \myifu/myicache/_1834_ ;
wire \myifu/myicache/_1835_ ;
wire \myifu/myicache/_1836_ ;
wire \myifu/myicache/_1837_ ;
wire \myifu/myicache/_1838_ ;
wire \myifu/myicache/_1839_ ;
wire \myifu/myicache/_1840_ ;
wire \myifu/myicache/_1841_ ;
wire \myifu/myicache/_1842_ ;
wire \myifu/myicache/_1843_ ;
wire \myifu/myicache/_1844_ ;
wire \myifu/myicache/_1845_ ;
wire \myifu/myicache/_1846_ ;
wire \myifu/myicache/_1847_ ;
wire \myifu/myicache/_1848_ ;
wire \myifu/myicache/_1849_ ;
wire \myifu/myicache/_1850_ ;
wire \myifu/myicache/_1851_ ;
wire \myifu/myicache/_1852_ ;
wire \myifu/myicache/_1853_ ;
wire \myifu/myicache/_1854_ ;
wire \myifu/myicache/_1855_ ;
wire \myifu/myicache/_1856_ ;
wire \myifu/myicache/_1857_ ;
wire \myifu/myicache/_1858_ ;
wire \myifu/myicache/_1859_ ;
wire \myifu/myicache/_1860_ ;
wire \myifu/myicache/_1861_ ;
wire \myifu/myicache/_1862_ ;
wire \myifu/myicache/_1863_ ;
wire \myifu/myicache/_1864_ ;
wire \myifu/myicache/_1865_ ;
wire \myifu/myicache/_1866_ ;
wire \myifu/myicache/_1867_ ;
wire \myifu/myicache/_1868_ ;
wire \myifu/myicache/_1869_ ;
wire \myifu/myicache/_1870_ ;
wire \myifu/myicache/_1871_ ;
wire \myifu/myicache/_1872_ ;
wire \myifu/myicache/_1873_ ;
wire \myifu/myicache/_1874_ ;
wire \myifu/myicache/_1875_ ;
wire \myifu/myicache/_1876_ ;
wire \myifu/myicache/_1877_ ;
wire \myifu/myicache/_1878_ ;
wire \myifu/myicache/_1879_ ;
wire \myifu/myicache/_1880_ ;
wire \myifu/myicache/_1881_ ;
wire \myifu/myicache/_1882_ ;
wire \myifu/myicache/_1883_ ;
wire \myifu/myicache/_1884_ ;
wire \myifu/myicache/_1885_ ;
wire \myifu/myicache/_1886_ ;
wire \myifu/myicache/_1887_ ;
wire \myifu/myicache/_1888_ ;
wire \myifu/myicache/_1889_ ;
wire \myifu/myicache/_1890_ ;
wire \myifu/myicache/_1891_ ;
wire \myifu/myicache/_1892_ ;
wire \myifu/myicache/_1893_ ;
wire \myifu/myicache/_1894_ ;
wire \myifu/myicache/_1895_ ;
wire \myifu/myicache/_1896_ ;
wire \myifu/myicache/_1897_ ;
wire \myifu/myicache/_1898_ ;
wire \myifu/myicache/_1899_ ;
wire \myifu/myicache/_1900_ ;
wire \myifu/myicache/_1901_ ;
wire \myifu/myicache/_1902_ ;
wire \myifu/myicache/_1903_ ;
wire \myifu/myicache/_1904_ ;
wire \myifu/myicache/_1905_ ;
wire \myifu/myicache/_1906_ ;
wire \myifu/myicache/_1907_ ;
wire \myifu/myicache/_1908_ ;
wire \myifu/myicache/_1909_ ;
wire \myifu/myicache/_1910_ ;
wire \myifu/myicache/_1911_ ;
wire \myifu/myicache/_1912_ ;
wire \myifu/myicache/_1913_ ;
wire \myifu/myicache/_1914_ ;
wire \myifu/myicache/_1915_ ;
wire \myifu/myicache/_1916_ ;
wire \myifu/myicache/_1917_ ;
wire \myifu/myicache/_1918_ ;
wire \myifu/myicache/_1919_ ;
wire \myifu/myicache/_1920_ ;
wire \myifu/myicache/_1921_ ;
wire \myifu/myicache/_1922_ ;
wire \myifu/myicache/_1923_ ;
wire \myifu/myicache/_1924_ ;
wire \myifu/myicache/_1925_ ;
wire \myifu/myicache/_1926_ ;
wire \myifu/myicache/_1927_ ;
wire \myifu/myicache/_1928_ ;
wire \myifu/myicache/_1929_ ;
wire \myifu/myicache/_1930_ ;
wire \myifu/myicache/_1931_ ;
wire \myifu/myicache/_1932_ ;
wire \myifu/myicache/_1933_ ;
wire \myifu/myicache/_1934_ ;
wire \myifu/myicache/_1935_ ;
wire \myifu/myicache/_1936_ ;
wire \myifu/myicache/_1937_ ;
wire \myifu/myicache/_1938_ ;
wire \myifu/myicache/_1939_ ;
wire \myifu/myicache/_1940_ ;
wire \myifu/myicache/_1941_ ;
wire \myifu/myicache/_1942_ ;
wire \myifu/myicache/_1943_ ;
wire \myifu/myicache/_1944_ ;
wire \myifu/myicache/_1945_ ;
wire \myifu/myicache/_1946_ ;
wire \myifu/myicache/_1947_ ;
wire \myifu/myicache/_1948_ ;
wire \myifu/myicache/_1949_ ;
wire \myifu/myicache/_1950_ ;
wire \myifu/myicache/_1951_ ;
wire \myifu/myicache/_1952_ ;
wire \myifu/myicache/_1953_ ;
wire \myifu/myicache/_1954_ ;
wire \myifu/myicache/_1955_ ;
wire \myifu/myicache/_1956_ ;
wire \myifu/myicache/_1957_ ;
wire \myifu/myicache/_1958_ ;
wire \myifu/myicache/_1959_ ;
wire \myifu/myicache/_1960_ ;
wire \myifu/myicache/_1961_ ;
wire \myifu/myicache/_1962_ ;
wire \myifu/myicache/_1963_ ;
wire \myifu/myicache/_1964_ ;
wire \myifu/myicache/_1965_ ;
wire \myifu/myicache/_1966_ ;
wire \myifu/myicache/_1967_ ;
wire \myifu/myicache/_1968_ ;
wire \myifu/myicache/_1969_ ;
wire \myifu/myicache/data[0][0] ;
wire \myifu/myicache/data[0][10] ;
wire \myifu/myicache/data[0][11] ;
wire \myifu/myicache/data[0][12] ;
wire \myifu/myicache/data[0][13] ;
wire \myifu/myicache/data[0][14] ;
wire \myifu/myicache/data[0][15] ;
wire \myifu/myicache/data[0][16] ;
wire \myifu/myicache/data[0][17] ;
wire \myifu/myicache/data[0][18] ;
wire \myifu/myicache/data[0][19] ;
wire \myifu/myicache/data[0][1] ;
wire \myifu/myicache/data[0][20] ;
wire \myifu/myicache/data[0][21] ;
wire \myifu/myicache/data[0][22] ;
wire \myifu/myicache/data[0][23] ;
wire \myifu/myicache/data[0][24] ;
wire \myifu/myicache/data[0][25] ;
wire \myifu/myicache/data[0][26] ;
wire \myifu/myicache/data[0][27] ;
wire \myifu/myicache/data[0][28] ;
wire \myifu/myicache/data[0][29] ;
wire \myifu/myicache/data[0][2] ;
wire \myifu/myicache/data[0][30] ;
wire \myifu/myicache/data[0][31] ;
wire \myifu/myicache/data[0][3] ;
wire \myifu/myicache/data[0][4] ;
wire \myifu/myicache/data[0][5] ;
wire \myifu/myicache/data[0][6] ;
wire \myifu/myicache/data[0][7] ;
wire \myifu/myicache/data[0][8] ;
wire \myifu/myicache/data[0][9] ;
wire \myifu/myicache/data[1][0] ;
wire \myifu/myicache/data[1][10] ;
wire \myifu/myicache/data[1][11] ;
wire \myifu/myicache/data[1][12] ;
wire \myifu/myicache/data[1][13] ;
wire \myifu/myicache/data[1][14] ;
wire \myifu/myicache/data[1][15] ;
wire \myifu/myicache/data[1][16] ;
wire \myifu/myicache/data[1][17] ;
wire \myifu/myicache/data[1][18] ;
wire \myifu/myicache/data[1][19] ;
wire \myifu/myicache/data[1][1] ;
wire \myifu/myicache/data[1][20] ;
wire \myifu/myicache/data[1][21] ;
wire \myifu/myicache/data[1][22] ;
wire \myifu/myicache/data[1][23] ;
wire \myifu/myicache/data[1][24] ;
wire \myifu/myicache/data[1][25] ;
wire \myifu/myicache/data[1][26] ;
wire \myifu/myicache/data[1][27] ;
wire \myifu/myicache/data[1][28] ;
wire \myifu/myicache/data[1][29] ;
wire \myifu/myicache/data[1][2] ;
wire \myifu/myicache/data[1][30] ;
wire \myifu/myicache/data[1][31] ;
wire \myifu/myicache/data[1][3] ;
wire \myifu/myicache/data[1][4] ;
wire \myifu/myicache/data[1][5] ;
wire \myifu/myicache/data[1][6] ;
wire \myifu/myicache/data[1][7] ;
wire \myifu/myicache/data[1][8] ;
wire \myifu/myicache/data[1][9] ;
wire \myifu/myicache/data[2][0] ;
wire \myifu/myicache/data[2][10] ;
wire \myifu/myicache/data[2][11] ;
wire \myifu/myicache/data[2][12] ;
wire \myifu/myicache/data[2][13] ;
wire \myifu/myicache/data[2][14] ;
wire \myifu/myicache/data[2][15] ;
wire \myifu/myicache/data[2][16] ;
wire \myifu/myicache/data[2][17] ;
wire \myifu/myicache/data[2][18] ;
wire \myifu/myicache/data[2][19] ;
wire \myifu/myicache/data[2][1] ;
wire \myifu/myicache/data[2][20] ;
wire \myifu/myicache/data[2][21] ;
wire \myifu/myicache/data[2][22] ;
wire \myifu/myicache/data[2][23] ;
wire \myifu/myicache/data[2][24] ;
wire \myifu/myicache/data[2][25] ;
wire \myifu/myicache/data[2][26] ;
wire \myifu/myicache/data[2][27] ;
wire \myifu/myicache/data[2][28] ;
wire \myifu/myicache/data[2][29] ;
wire \myifu/myicache/data[2][2] ;
wire \myifu/myicache/data[2][30] ;
wire \myifu/myicache/data[2][31] ;
wire \myifu/myicache/data[2][3] ;
wire \myifu/myicache/data[2][4] ;
wire \myifu/myicache/data[2][5] ;
wire \myifu/myicache/data[2][6] ;
wire \myifu/myicache/data[2][7] ;
wire \myifu/myicache/data[2][8] ;
wire \myifu/myicache/data[2][9] ;
wire \myifu/myicache/data[3][0] ;
wire \myifu/myicache/data[3][10] ;
wire \myifu/myicache/data[3][11] ;
wire \myifu/myicache/data[3][12] ;
wire \myifu/myicache/data[3][13] ;
wire \myifu/myicache/data[3][14] ;
wire \myifu/myicache/data[3][15] ;
wire \myifu/myicache/data[3][16] ;
wire \myifu/myicache/data[3][17] ;
wire \myifu/myicache/data[3][18] ;
wire \myifu/myicache/data[3][19] ;
wire \myifu/myicache/data[3][1] ;
wire \myifu/myicache/data[3][20] ;
wire \myifu/myicache/data[3][21] ;
wire \myifu/myicache/data[3][22] ;
wire \myifu/myicache/data[3][23] ;
wire \myifu/myicache/data[3][24] ;
wire \myifu/myicache/data[3][25] ;
wire \myifu/myicache/data[3][26] ;
wire \myifu/myicache/data[3][27] ;
wire \myifu/myicache/data[3][28] ;
wire \myifu/myicache/data[3][29] ;
wire \myifu/myicache/data[3][2] ;
wire \myifu/myicache/data[3][30] ;
wire \myifu/myicache/data[3][31] ;
wire \myifu/myicache/data[3][3] ;
wire \myifu/myicache/data[3][4] ;
wire \myifu/myicache/data[3][5] ;
wire \myifu/myicache/data[3][6] ;
wire \myifu/myicache/data[3][7] ;
wire \myifu/myicache/data[3][8] ;
wire \myifu/myicache/data[3][9] ;
wire \myifu/myicache/data[4][0] ;
wire \myifu/myicache/data[4][10] ;
wire \myifu/myicache/data[4][11] ;
wire \myifu/myicache/data[4][12] ;
wire \myifu/myicache/data[4][13] ;
wire \myifu/myicache/data[4][14] ;
wire \myifu/myicache/data[4][15] ;
wire \myifu/myicache/data[4][16] ;
wire \myifu/myicache/data[4][17] ;
wire \myifu/myicache/data[4][18] ;
wire \myifu/myicache/data[4][19] ;
wire \myifu/myicache/data[4][1] ;
wire \myifu/myicache/data[4][20] ;
wire \myifu/myicache/data[4][21] ;
wire \myifu/myicache/data[4][22] ;
wire \myifu/myicache/data[4][23] ;
wire \myifu/myicache/data[4][24] ;
wire \myifu/myicache/data[4][25] ;
wire \myifu/myicache/data[4][26] ;
wire \myifu/myicache/data[4][27] ;
wire \myifu/myicache/data[4][28] ;
wire \myifu/myicache/data[4][29] ;
wire \myifu/myicache/data[4][2] ;
wire \myifu/myicache/data[4][30] ;
wire \myifu/myicache/data[4][31] ;
wire \myifu/myicache/data[4][3] ;
wire \myifu/myicache/data[4][4] ;
wire \myifu/myicache/data[4][5] ;
wire \myifu/myicache/data[4][6] ;
wire \myifu/myicache/data[4][7] ;
wire \myifu/myicache/data[4][8] ;
wire \myifu/myicache/data[4][9] ;
wire \myifu/myicache/data[5][0] ;
wire \myifu/myicache/data[5][10] ;
wire \myifu/myicache/data[5][11] ;
wire \myifu/myicache/data[5][12] ;
wire \myifu/myicache/data[5][13] ;
wire \myifu/myicache/data[5][14] ;
wire \myifu/myicache/data[5][15] ;
wire \myifu/myicache/data[5][16] ;
wire \myifu/myicache/data[5][17] ;
wire \myifu/myicache/data[5][18] ;
wire \myifu/myicache/data[5][19] ;
wire \myifu/myicache/data[5][1] ;
wire \myifu/myicache/data[5][20] ;
wire \myifu/myicache/data[5][21] ;
wire \myifu/myicache/data[5][22] ;
wire \myifu/myicache/data[5][23] ;
wire \myifu/myicache/data[5][24] ;
wire \myifu/myicache/data[5][25] ;
wire \myifu/myicache/data[5][26] ;
wire \myifu/myicache/data[5][27] ;
wire \myifu/myicache/data[5][28] ;
wire \myifu/myicache/data[5][29] ;
wire \myifu/myicache/data[5][2] ;
wire \myifu/myicache/data[5][30] ;
wire \myifu/myicache/data[5][31] ;
wire \myifu/myicache/data[5][3] ;
wire \myifu/myicache/data[5][4] ;
wire \myifu/myicache/data[5][5] ;
wire \myifu/myicache/data[5][6] ;
wire \myifu/myicache/data[5][7] ;
wire \myifu/myicache/data[5][8] ;
wire \myifu/myicache/data[5][9] ;
wire \myifu/myicache/data[6][0] ;
wire \myifu/myicache/data[6][10] ;
wire \myifu/myicache/data[6][11] ;
wire \myifu/myicache/data[6][12] ;
wire \myifu/myicache/data[6][13] ;
wire \myifu/myicache/data[6][14] ;
wire \myifu/myicache/data[6][15] ;
wire \myifu/myicache/data[6][16] ;
wire \myifu/myicache/data[6][17] ;
wire \myifu/myicache/data[6][18] ;
wire \myifu/myicache/data[6][19] ;
wire \myifu/myicache/data[6][1] ;
wire \myifu/myicache/data[6][20] ;
wire \myifu/myicache/data[6][21] ;
wire \myifu/myicache/data[6][22] ;
wire \myifu/myicache/data[6][23] ;
wire \myifu/myicache/data[6][24] ;
wire \myifu/myicache/data[6][25] ;
wire \myifu/myicache/data[6][26] ;
wire \myifu/myicache/data[6][27] ;
wire \myifu/myicache/data[6][28] ;
wire \myifu/myicache/data[6][29] ;
wire \myifu/myicache/data[6][2] ;
wire \myifu/myicache/data[6][30] ;
wire \myifu/myicache/data[6][31] ;
wire \myifu/myicache/data[6][3] ;
wire \myifu/myicache/data[6][4] ;
wire \myifu/myicache/data[6][5] ;
wire \myifu/myicache/data[6][6] ;
wire \myifu/myicache/data[6][7] ;
wire \myifu/myicache/data[6][8] ;
wire \myifu/myicache/data[6][9] ;
wire \myifu/myicache/data[7][0] ;
wire \myifu/myicache/data[7][10] ;
wire \myifu/myicache/data[7][11] ;
wire \myifu/myicache/data[7][12] ;
wire \myifu/myicache/data[7][13] ;
wire \myifu/myicache/data[7][14] ;
wire \myifu/myicache/data[7][15] ;
wire \myifu/myicache/data[7][16] ;
wire \myifu/myicache/data[7][17] ;
wire \myifu/myicache/data[7][18] ;
wire \myifu/myicache/data[7][19] ;
wire \myifu/myicache/data[7][1] ;
wire \myifu/myicache/data[7][20] ;
wire \myifu/myicache/data[7][21] ;
wire \myifu/myicache/data[7][22] ;
wire \myifu/myicache/data[7][23] ;
wire \myifu/myicache/data[7][24] ;
wire \myifu/myicache/data[7][25] ;
wire \myifu/myicache/data[7][26] ;
wire \myifu/myicache/data[7][27] ;
wire \myifu/myicache/data[7][28] ;
wire \myifu/myicache/data[7][29] ;
wire \myifu/myicache/data[7][2] ;
wire \myifu/myicache/data[7][30] ;
wire \myifu/myicache/data[7][31] ;
wire \myifu/myicache/data[7][3] ;
wire \myifu/myicache/data[7][4] ;
wire \myifu/myicache/data[7][5] ;
wire \myifu/myicache/data[7][6] ;
wire \myifu/myicache/data[7][7] ;
wire \myifu/myicache/data[7][8] ;
wire \myifu/myicache/data[7][9] ;
wire \myifu/myicache/tag[0][0] ;
wire \myifu/myicache/tag[0][10] ;
wire \myifu/myicache/tag[0][11] ;
wire \myifu/myicache/tag[0][12] ;
wire \myifu/myicache/tag[0][13] ;
wire \myifu/myicache/tag[0][14] ;
wire \myifu/myicache/tag[0][15] ;
wire \myifu/myicache/tag[0][16] ;
wire \myifu/myicache/tag[0][17] ;
wire \myifu/myicache/tag[0][18] ;
wire \myifu/myicache/tag[0][19] ;
wire \myifu/myicache/tag[0][1] ;
wire \myifu/myicache/tag[0][20] ;
wire \myifu/myicache/tag[0][21] ;
wire \myifu/myicache/tag[0][22] ;
wire \myifu/myicache/tag[0][23] ;
wire \myifu/myicache/tag[0][24] ;
wire \myifu/myicache/tag[0][25] ;
wire \myifu/myicache/tag[0][26] ;
wire \myifu/myicache/tag[0][2] ;
wire \myifu/myicache/tag[0][3] ;
wire \myifu/myicache/tag[0][4] ;
wire \myifu/myicache/tag[0][5] ;
wire \myifu/myicache/tag[0][6] ;
wire \myifu/myicache/tag[0][7] ;
wire \myifu/myicache/tag[0][8] ;
wire \myifu/myicache/tag[0][9] ;
wire \myifu/myicache/tag[1][0] ;
wire \myifu/myicache/tag[1][10] ;
wire \myifu/myicache/tag[1][11] ;
wire \myifu/myicache/tag[1][12] ;
wire \myifu/myicache/tag[1][13] ;
wire \myifu/myicache/tag[1][14] ;
wire \myifu/myicache/tag[1][15] ;
wire \myifu/myicache/tag[1][16] ;
wire \myifu/myicache/tag[1][17] ;
wire \myifu/myicache/tag[1][18] ;
wire \myifu/myicache/tag[1][19] ;
wire \myifu/myicache/tag[1][1] ;
wire \myifu/myicache/tag[1][20] ;
wire \myifu/myicache/tag[1][21] ;
wire \myifu/myicache/tag[1][22] ;
wire \myifu/myicache/tag[1][23] ;
wire \myifu/myicache/tag[1][24] ;
wire \myifu/myicache/tag[1][25] ;
wire \myifu/myicache/tag[1][26] ;
wire \myifu/myicache/tag[1][2] ;
wire \myifu/myicache/tag[1][3] ;
wire \myifu/myicache/tag[1][4] ;
wire \myifu/myicache/tag[1][5] ;
wire \myifu/myicache/tag[1][6] ;
wire \myifu/myicache/tag[1][7] ;
wire \myifu/myicache/tag[1][8] ;
wire \myifu/myicache/tag[1][9] ;
wire \myifu/myicache/tag[2][0] ;
wire \myifu/myicache/tag[2][10] ;
wire \myifu/myicache/tag[2][11] ;
wire \myifu/myicache/tag[2][12] ;
wire \myifu/myicache/tag[2][13] ;
wire \myifu/myicache/tag[2][14] ;
wire \myifu/myicache/tag[2][15] ;
wire \myifu/myicache/tag[2][16] ;
wire \myifu/myicache/tag[2][17] ;
wire \myifu/myicache/tag[2][18] ;
wire \myifu/myicache/tag[2][19] ;
wire \myifu/myicache/tag[2][1] ;
wire \myifu/myicache/tag[2][20] ;
wire \myifu/myicache/tag[2][21] ;
wire \myifu/myicache/tag[2][22] ;
wire \myifu/myicache/tag[2][23] ;
wire \myifu/myicache/tag[2][24] ;
wire \myifu/myicache/tag[2][25] ;
wire \myifu/myicache/tag[2][26] ;
wire \myifu/myicache/tag[2][2] ;
wire \myifu/myicache/tag[2][3] ;
wire \myifu/myicache/tag[2][4] ;
wire \myifu/myicache/tag[2][5] ;
wire \myifu/myicache/tag[2][6] ;
wire \myifu/myicache/tag[2][7] ;
wire \myifu/myicache/tag[2][8] ;
wire \myifu/myicache/tag[2][9] ;
wire \myifu/myicache/tag[3][0] ;
wire \myifu/myicache/tag[3][10] ;
wire \myifu/myicache/tag[3][11] ;
wire \myifu/myicache/tag[3][12] ;
wire \myifu/myicache/tag[3][13] ;
wire \myifu/myicache/tag[3][14] ;
wire \myifu/myicache/tag[3][15] ;
wire \myifu/myicache/tag[3][16] ;
wire \myifu/myicache/tag[3][17] ;
wire \myifu/myicache/tag[3][18] ;
wire \myifu/myicache/tag[3][19] ;
wire \myifu/myicache/tag[3][1] ;
wire \myifu/myicache/tag[3][20] ;
wire \myifu/myicache/tag[3][21] ;
wire \myifu/myicache/tag[3][22] ;
wire \myifu/myicache/tag[3][23] ;
wire \myifu/myicache/tag[3][24] ;
wire \myifu/myicache/tag[3][25] ;
wire \myifu/myicache/tag[3][26] ;
wire \myifu/myicache/tag[3][2] ;
wire \myifu/myicache/tag[3][3] ;
wire \myifu/myicache/tag[3][4] ;
wire \myifu/myicache/tag[3][5] ;
wire \myifu/myicache/tag[3][6] ;
wire \myifu/myicache/tag[3][7] ;
wire \myifu/myicache/tag[3][8] ;
wire \myifu/myicache/tag[3][9] ;
wire \mylsu/_0000_ ;
wire \mylsu/_0001_ ;
wire \mylsu/_0002_ ;
wire \mylsu/_0003_ ;
wire \mylsu/_0004_ ;
wire \mylsu/_0005_ ;
wire \mylsu/_0006_ ;
wire \mylsu/_0007_ ;
wire \mylsu/_0008_ ;
wire \mylsu/_0009_ ;
wire \mylsu/_0010_ ;
wire \mylsu/_0011_ ;
wire \mylsu/_0012_ ;
wire \mylsu/_0013_ ;
wire \mylsu/_0014_ ;
wire \mylsu/_0015_ ;
wire \mylsu/_0016_ ;
wire \mylsu/_0017_ ;
wire \mylsu/_0018_ ;
wire \mylsu/_0019_ ;
wire \mylsu/_0020_ ;
wire \mylsu/_0021_ ;
wire \mylsu/_0022_ ;
wire \mylsu/_0023_ ;
wire \mylsu/_0024_ ;
wire \mylsu/_0025_ ;
wire \mylsu/_0026_ ;
wire \mylsu/_0027_ ;
wire \mylsu/_0028_ ;
wire \mylsu/_0029_ ;
wire \mylsu/_0030_ ;
wire \mylsu/_0031_ ;
wire \mylsu/_0032_ ;
wire \mylsu/_0033_ ;
wire \mylsu/_0034_ ;
wire \mylsu/_0035_ ;
wire \mylsu/_0036_ ;
wire \mylsu/_0037_ ;
wire \mylsu/_0038_ ;
wire \mylsu/_0039_ ;
wire \mylsu/_0040_ ;
wire \mylsu/_0041_ ;
wire \mylsu/_0042_ ;
wire \mylsu/_0043_ ;
wire \mylsu/_0044_ ;
wire \mylsu/_0045_ ;
wire \mylsu/_0046_ ;
wire \mylsu/_0047_ ;
wire \mylsu/_0048_ ;
wire \mylsu/_0049_ ;
wire \mylsu/_0050_ ;
wire \mylsu/_0051_ ;
wire \mylsu/_0052_ ;
wire \mylsu/_0053_ ;
wire \mylsu/_0054_ ;
wire \mylsu/_0055_ ;
wire \mylsu/_0056_ ;
wire \mylsu/_0057_ ;
wire \mylsu/_0058_ ;
wire \mylsu/_0059_ ;
wire \mylsu/_0060_ ;
wire \mylsu/_0061_ ;
wire \mylsu/_0062_ ;
wire \mylsu/_0063_ ;
wire \mylsu/_0064_ ;
wire \mylsu/_0065_ ;
wire \mylsu/_0066_ ;
wire \mylsu/_0067_ ;
wire \mylsu/_0068_ ;
wire \mylsu/_0069_ ;
wire \mylsu/_0070_ ;
wire \mylsu/_0071_ ;
wire \mylsu/_0072_ ;
wire \mylsu/_0073_ ;
wire \mylsu/_0074_ ;
wire \mylsu/_0075_ ;
wire \mylsu/_0076_ ;
wire \mylsu/_0077_ ;
wire \mylsu/_0078_ ;
wire \mylsu/_0079_ ;
wire \mylsu/_0080_ ;
wire \mylsu/_0081_ ;
wire \mylsu/_0082_ ;
wire \mylsu/_0083_ ;
wire \mylsu/_0084_ ;
wire \mylsu/_0085_ ;
wire \mylsu/_0086_ ;
wire \mylsu/_0087_ ;
wire \mylsu/_0088_ ;
wire \mylsu/_0089_ ;
wire \mylsu/_0090_ ;
wire \mylsu/_0091_ ;
wire \mylsu/_0092_ ;
wire \mylsu/_0093_ ;
wire \mylsu/_0094_ ;
wire \mylsu/_0095_ ;
wire \mylsu/_0096_ ;
wire \mylsu/_0097_ ;
wire \mylsu/_0098_ ;
wire \mylsu/_0099_ ;
wire \mylsu/_0100_ ;
wire \mylsu/_0101_ ;
wire \mylsu/_0102_ ;
wire \mylsu/_0103_ ;
wire \mylsu/_0104_ ;
wire \mylsu/_0105_ ;
wire \mylsu/_0106_ ;
wire \mylsu/_0107_ ;
wire \mylsu/_0108_ ;
wire \mylsu/_0109_ ;
wire \mylsu/_0110_ ;
wire \mylsu/_0111_ ;
wire \mylsu/_0112_ ;
wire \mylsu/_0113_ ;
wire \mylsu/_0114_ ;
wire \mylsu/_0115_ ;
wire \mylsu/_0116_ ;
wire \mylsu/_0117_ ;
wire \mylsu/_0118_ ;
wire \mylsu/_0119_ ;
wire \mylsu/_0120_ ;
wire \mylsu/_0121_ ;
wire \mylsu/_0122_ ;
wire \mylsu/_0123_ ;
wire \mylsu/_0124_ ;
wire \mylsu/_0125_ ;
wire \mylsu/_0126_ ;
wire \mylsu/_0127_ ;
wire \mylsu/_0128_ ;
wire \mylsu/_0129_ ;
wire \mylsu/_0130_ ;
wire \mylsu/_0131_ ;
wire \mylsu/_0132_ ;
wire \mylsu/_0133_ ;
wire \mylsu/_0134_ ;
wire \mylsu/_0135_ ;
wire \mylsu/_0136_ ;
wire \mylsu/_0137_ ;
wire \mylsu/_0138_ ;
wire \mylsu/_0139_ ;
wire \mylsu/_0140_ ;
wire \mylsu/_0141_ ;
wire \mylsu/_0142_ ;
wire \mylsu/_0143_ ;
wire \mylsu/_0144_ ;
wire \mylsu/_0145_ ;
wire \mylsu/_0146_ ;
wire \mylsu/_0147_ ;
wire \mylsu/_0148_ ;
wire \mylsu/_0149_ ;
wire \mylsu/_0150_ ;
wire \mylsu/_0151_ ;
wire \mylsu/_0152_ ;
wire \mylsu/_0153_ ;
wire \mylsu/_0154_ ;
wire \mylsu/_0155_ ;
wire \mylsu/_0156_ ;
wire \mylsu/_0157_ ;
wire \mylsu/_0158_ ;
wire \mylsu/_0159_ ;
wire \mylsu/_0160_ ;
wire \mylsu/_0161_ ;
wire \mylsu/_0162_ ;
wire \mylsu/_0163_ ;
wire \mylsu/_0164_ ;
wire \mylsu/_0165_ ;
wire \mylsu/_0166_ ;
wire \mylsu/_0167_ ;
wire \mylsu/_0168_ ;
wire \mylsu/_0169_ ;
wire \mylsu/_0170_ ;
wire \mylsu/_0171_ ;
wire \mylsu/_0172_ ;
wire \mylsu/_0173_ ;
wire \mylsu/_0174_ ;
wire \mylsu/_0175_ ;
wire \mylsu/_0176_ ;
wire \mylsu/_0177_ ;
wire \mylsu/_0178_ ;
wire \mylsu/_0179_ ;
wire \mylsu/_0180_ ;
wire \mylsu/_0181_ ;
wire \mylsu/_0182_ ;
wire \mylsu/_0183_ ;
wire \mylsu/_0184_ ;
wire \mylsu/_0185_ ;
wire \mylsu/_0186_ ;
wire \mylsu/_0187_ ;
wire \mylsu/_0188_ ;
wire \mylsu/_0189_ ;
wire \mylsu/_0190_ ;
wire \mylsu/_0191_ ;
wire \mylsu/_0192_ ;
wire \mylsu/_0193_ ;
wire \mylsu/_0194_ ;
wire \mylsu/_0195_ ;
wire \mylsu/_0196_ ;
wire \mylsu/_0197_ ;
wire \mylsu/_0198_ ;
wire \mylsu/_0199_ ;
wire \mylsu/_0200_ ;
wire \mylsu/_0201_ ;
wire \mylsu/_0202_ ;
wire \mylsu/_0203_ ;
wire \mylsu/_0204_ ;
wire \mylsu/_0205_ ;
wire \mylsu/_0206_ ;
wire \mylsu/_0207_ ;
wire \mylsu/_0208_ ;
wire \mylsu/_0209_ ;
wire \mylsu/_0210_ ;
wire \mylsu/_0211_ ;
wire \mylsu/_0212_ ;
wire \mylsu/_0213_ ;
wire \mylsu/_0214_ ;
wire \mylsu/_0215_ ;
wire \mylsu/_0216_ ;
wire \mylsu/_0217_ ;
wire \mylsu/_0218_ ;
wire \mylsu/_0219_ ;
wire \mylsu/_0220_ ;
wire \mylsu/_0221_ ;
wire \mylsu/_0222_ ;
wire \mylsu/_0223_ ;
wire \mylsu/_0224_ ;
wire \mylsu/_0225_ ;
wire \mylsu/_0226_ ;
wire \mylsu/_0227_ ;
wire \mylsu/_0228_ ;
wire \mylsu/_0229_ ;
wire \mylsu/_0230_ ;
wire \mylsu/_0231_ ;
wire \mylsu/_0232_ ;
wire \mylsu/_0233_ ;
wire \mylsu/_0234_ ;
wire \mylsu/_0235_ ;
wire \mylsu/_0236_ ;
wire \mylsu/_0237_ ;
wire \mylsu/_0238_ ;
wire \mylsu/_0239_ ;
wire \mylsu/_0240_ ;
wire \mylsu/_0241_ ;
wire \mylsu/_0242_ ;
wire \mylsu/_0243_ ;
wire \mylsu/_0244_ ;
wire \mylsu/_0245_ ;
wire \mylsu/_0246_ ;
wire \mylsu/_0247_ ;
wire \mylsu/_0248_ ;
wire \mylsu/_0249_ ;
wire \mylsu/_0250_ ;
wire \mylsu/_0251_ ;
wire \mylsu/_0252_ ;
wire \mylsu/_0253_ ;
wire \mylsu/_0254_ ;
wire \mylsu/_0255_ ;
wire \mylsu/_0256_ ;
wire \mylsu/_0257_ ;
wire \mylsu/_0258_ ;
wire \mylsu/_0259_ ;
wire \mylsu/_0260_ ;
wire \mylsu/_0261_ ;
wire \mylsu/_0262_ ;
wire \mylsu/_0263_ ;
wire \mylsu/_0264_ ;
wire \mylsu/_0265_ ;
wire \mylsu/_0266_ ;
wire \mylsu/_0267_ ;
wire \mylsu/_0268_ ;
wire \mylsu/_0269_ ;
wire \mylsu/_0270_ ;
wire \mylsu/_0271_ ;
wire \mylsu/_0272_ ;
wire \mylsu/_0273_ ;
wire \mylsu/_0274_ ;
wire \mylsu/_0275_ ;
wire \mylsu/_0276_ ;
wire \mylsu/_0277_ ;
wire \mylsu/_0278_ ;
wire \mylsu/_0279_ ;
wire \mylsu/_0280_ ;
wire \mylsu/_0281_ ;
wire \mylsu/_0282_ ;
wire \mylsu/_0283_ ;
wire \mylsu/_0284_ ;
wire \mylsu/_0285_ ;
wire \mylsu/_0286_ ;
wire \mylsu/_0287_ ;
wire \mylsu/_0288_ ;
wire \mylsu/_0289_ ;
wire \mylsu/_0290_ ;
wire \mylsu/_0291_ ;
wire \mylsu/_0292_ ;
wire \mylsu/_0293_ ;
wire \mylsu/_0294_ ;
wire \mylsu/_0295_ ;
wire \mylsu/_0296_ ;
wire \mylsu/_0297_ ;
wire \mylsu/_0298_ ;
wire \mylsu/_0299_ ;
wire \mylsu/_0300_ ;
wire \mylsu/_0301_ ;
wire \mylsu/_0302_ ;
wire \mylsu/_0303_ ;
wire \mylsu/_0304_ ;
wire \mylsu/_0305_ ;
wire \mylsu/_0306_ ;
wire \mylsu/_0307_ ;
wire \mylsu/_0308_ ;
wire \mylsu/_0309_ ;
wire \mylsu/_0310_ ;
wire \mylsu/_0311_ ;
wire \mylsu/_0312_ ;
wire \mylsu/_0313_ ;
wire \mylsu/_0314_ ;
wire \mylsu/_0315_ ;
wire \mylsu/_0316_ ;
wire \mylsu/_0317_ ;
wire \mylsu/_0318_ ;
wire \mylsu/_0319_ ;
wire \mylsu/_0320_ ;
wire \mylsu/_0321_ ;
wire \mylsu/_0322_ ;
wire \mylsu/_0323_ ;
wire \mylsu/_0324_ ;
wire \mylsu/_0325_ ;
wire \mylsu/_0326_ ;
wire \mylsu/_0327_ ;
wire \mylsu/_0328_ ;
wire \mylsu/_0329_ ;
wire \mylsu/_0330_ ;
wire \mylsu/_0331_ ;
wire \mylsu/_0332_ ;
wire \mylsu/_0333_ ;
wire \mylsu/_0334_ ;
wire \mylsu/_0335_ ;
wire \mylsu/_0336_ ;
wire \mylsu/_0337_ ;
wire \mylsu/_0338_ ;
wire \mylsu/_0339_ ;
wire \mylsu/_0340_ ;
wire \mylsu/_0341_ ;
wire \mylsu/_0342_ ;
wire \mylsu/_0343_ ;
wire \mylsu/_0344_ ;
wire \mylsu/_0345_ ;
wire \mylsu/_0346_ ;
wire \mylsu/_0347_ ;
wire \mylsu/_0348_ ;
wire \mylsu/_0349_ ;
wire \mylsu/_0350_ ;
wire \mylsu/_0351_ ;
wire \mylsu/_0352_ ;
wire \mylsu/_0353_ ;
wire \mylsu/_0354_ ;
wire \mylsu/_0355_ ;
wire \mylsu/_0356_ ;
wire \mylsu/_0357_ ;
wire \mylsu/_0358_ ;
wire \mylsu/_0359_ ;
wire \mylsu/_0360_ ;
wire \mylsu/_0361_ ;
wire \mylsu/_0362_ ;
wire \mylsu/_0363_ ;
wire \mylsu/_0364_ ;
wire \mylsu/_0365_ ;
wire \mylsu/_0366_ ;
wire \mylsu/_0367_ ;
wire \mylsu/_0368_ ;
wire \mylsu/_0369_ ;
wire \mylsu/_0370_ ;
wire \mylsu/_0371_ ;
wire \mylsu/_0372_ ;
wire \mylsu/_0373_ ;
wire \mylsu/_0374_ ;
wire \mylsu/_0375_ ;
wire \mylsu/_0376_ ;
wire \mylsu/_0377_ ;
wire \mylsu/_0378_ ;
wire \mylsu/_0379_ ;
wire \mylsu/_0380_ ;
wire \mylsu/_0381_ ;
wire \mylsu/_0382_ ;
wire \mylsu/_0383_ ;
wire \mylsu/_0384_ ;
wire \mylsu/_0385_ ;
wire \mylsu/_0386_ ;
wire \mylsu/_0387_ ;
wire \mylsu/_0388_ ;
wire \mylsu/_0389_ ;
wire \mylsu/_0390_ ;
wire \mylsu/_0391_ ;
wire \mylsu/_0392_ ;
wire \mylsu/_0393_ ;
wire \mylsu/_0394_ ;
wire \mylsu/_0395_ ;
wire \mylsu/_0396_ ;
wire \mylsu/_0397_ ;
wire \mylsu/_0398_ ;
wire \mylsu/_0399_ ;
wire \mylsu/_0400_ ;
wire \mylsu/_0401_ ;
wire \mylsu/_0402_ ;
wire \mylsu/_0403_ ;
wire \mylsu/_0404_ ;
wire \mylsu/_0405_ ;
wire \mylsu/_0406_ ;
wire \mylsu/_0407_ ;
wire \mylsu/_0408_ ;
wire \mylsu/_0409_ ;
wire \mylsu/_0410_ ;
wire \mylsu/_0411_ ;
wire \mylsu/_0412_ ;
wire \mylsu/_0413_ ;
wire \mylsu/_0414_ ;
wire \mylsu/_0415_ ;
wire \mylsu/_0416_ ;
wire \mylsu/_0417_ ;
wire \mylsu/_0418_ ;
wire \mylsu/_0419_ ;
wire \mylsu/_0420_ ;
wire \mylsu/_0421_ ;
wire \mylsu/_0422_ ;
wire \mylsu/_0423_ ;
wire \mylsu/_0424_ ;
wire \mylsu/_0425_ ;
wire \mylsu/_0426_ ;
wire \mylsu/_0427_ ;
wire \mylsu/_0428_ ;
wire \mylsu/_0429_ ;
wire \mylsu/_0430_ ;
wire \mylsu/_0431_ ;
wire \mylsu/_0432_ ;
wire \mylsu/_0433_ ;
wire \mylsu/_0434_ ;
wire \mylsu/_0435_ ;
wire \mylsu/_0436_ ;
wire \mylsu/_0437_ ;
wire \mylsu/_0438_ ;
wire \mylsu/_0439_ ;
wire \mylsu/_0440_ ;
wire \mylsu/_0441_ ;
wire \mylsu/_0442_ ;
wire \mylsu/_0443_ ;
wire \mylsu/_0444_ ;
wire \mylsu/_0445_ ;
wire \mylsu/_0446_ ;
wire \mylsu/_0447_ ;
wire \mylsu/_0448_ ;
wire \mylsu/_0449_ ;
wire \mylsu/_0450_ ;
wire \mylsu/_0451_ ;
wire \mylsu/_0452_ ;
wire \mylsu/_0453_ ;
wire \mylsu/_0454_ ;
wire \mylsu/_0455_ ;
wire \mylsu/_0456_ ;
wire \mylsu/_0457_ ;
wire \mylsu/_0458_ ;
wire \mylsu/_0459_ ;
wire \mylsu/_0460_ ;
wire \mylsu/_0461_ ;
wire \mylsu/_0462_ ;
wire \mylsu/_0463_ ;
wire \mylsu/_0464_ ;
wire \mylsu/_0465_ ;
wire \mylsu/_0466_ ;
wire \mylsu/_0467_ ;
wire \mylsu/_0468_ ;
wire \mylsu/_0469_ ;
wire \mylsu/_0470_ ;
wire \mylsu/_0471_ ;
wire \mylsu/_0472_ ;
wire \mylsu/_0473_ ;
wire \mylsu/_0474_ ;
wire \mylsu/_0475_ ;
wire \mylsu/_0476_ ;
wire \mylsu/_0477_ ;
wire \mylsu/_0478_ ;
wire \mylsu/_0479_ ;
wire \mylsu/_0480_ ;
wire \mylsu/_0481_ ;
wire \mylsu/_0482_ ;
wire \mylsu/_0483_ ;
wire \mylsu/_0484_ ;
wire \mylsu/_0485_ ;
wire \mylsu/_0486_ ;
wire \mylsu/_0487_ ;
wire \mylsu/_0488_ ;
wire \mylsu/_0489_ ;
wire \mylsu/_0490_ ;
wire \mylsu/_0491_ ;
wire \mylsu/_0492_ ;
wire \mylsu/_0493_ ;
wire \mylsu/_0494_ ;
wire \mylsu/_0495_ ;
wire \mylsu/_0496_ ;
wire \mylsu/_0497_ ;
wire \mylsu/_0498_ ;
wire \mylsu/_0499_ ;
wire \mylsu/_0500_ ;
wire \mylsu/_0501_ ;
wire \mylsu/_0502_ ;
wire \mylsu/_0503_ ;
wire \mylsu/_0504_ ;
wire \mylsu/_0505_ ;
wire \mylsu/_0506_ ;
wire \mylsu/_0507_ ;
wire \mylsu/_0508_ ;
wire \mylsu/_0509_ ;
wire \mylsu/_0510_ ;
wire \mylsu/_0511_ ;
wire \mylsu/_0512_ ;
wire \mylsu/_0513_ ;
wire \mylsu/_0514_ ;
wire \mylsu/_0515_ ;
wire \mylsu/_0516_ ;
wire \mylsu/_0517_ ;
wire \mylsu/_0518_ ;
wire \mylsu/_0519_ ;
wire \mylsu/_0520_ ;
wire \mylsu/_0521_ ;
wire \mylsu/_0522_ ;
wire \mylsu/_0523_ ;
wire \mylsu/_0524_ ;
wire \mylsu/_0525_ ;
wire \mylsu/_0526_ ;
wire \mylsu/_0527_ ;
wire \mylsu/_0528_ ;
wire \mylsu/_0529_ ;
wire \mylsu/_0530_ ;
wire \mylsu/_0531_ ;
wire \mylsu/_0532_ ;
wire \mylsu/_0533_ ;
wire \mylsu/_0534_ ;
wire \mylsu/_0535_ ;
wire \mylsu/_0536_ ;
wire \mylsu/_0537_ ;
wire \mylsu/_0538_ ;
wire \mylsu/_0539_ ;
wire \mylsu/_0540_ ;
wire \mylsu/_0541_ ;
wire \mylsu/_0542_ ;
wire \mylsu/_0543_ ;
wire \mylsu/_0544_ ;
wire \mylsu/_0545_ ;
wire \mylsu/_0546_ ;
wire \mylsu/_0547_ ;
wire \mylsu/_0548_ ;
wire \mylsu/_0549_ ;
wire \mylsu/_0550_ ;
wire \mylsu/_0551_ ;
wire \mylsu/_0552_ ;
wire \mylsu/_0553_ ;
wire \mylsu/_0554_ ;
wire \mylsu/_0555_ ;
wire \mylsu/_0556_ ;
wire \mylsu/_0557_ ;
wire \mylsu/_0558_ ;
wire \mylsu/_0559_ ;
wire \mylsu/_0560_ ;
wire \mylsu/_0561_ ;
wire \mylsu/_0562_ ;
wire \mylsu/_0563_ ;
wire \mylsu/_0564_ ;
wire \mylsu/_0565_ ;
wire \mylsu/_0566_ ;
wire \mylsu/_0567_ ;
wire \mylsu/_0568_ ;
wire \mylsu/_0569_ ;
wire \mylsu/_0570_ ;
wire \mylsu/_0571_ ;
wire \mylsu/_0572_ ;
wire \mylsu/_0573_ ;
wire \mylsu/_0574_ ;
wire \mylsu/_0575_ ;
wire \mylsu/_0576_ ;
wire \mylsu/_0577_ ;
wire \mylsu/_0578_ ;
wire \mylsu/_0579_ ;
wire \mylsu/_0580_ ;
wire \mylsu/_0581_ ;
wire \mylsu/_0582_ ;
wire \mylsu/_0583_ ;
wire \mylsu/_0584_ ;
wire \mylsu/_0585_ ;
wire \mylsu/_0586_ ;
wire \mylsu/_0587_ ;
wire \mylsu/_0588_ ;
wire \mylsu/_0589_ ;
wire \mylsu/_0590_ ;
wire \mylsu/_0591_ ;
wire \mylsu/_0592_ ;
wire \mylsu/_0593_ ;
wire \mylsu/_0594_ ;
wire \mylsu/_0595_ ;
wire \mylsu/_0596_ ;
wire \mylsu/_0597_ ;
wire \mylsu/_0598_ ;
wire \mylsu/_0599_ ;
wire \mylsu/_0600_ ;
wire \mylsu/_0601_ ;
wire \mylsu/_0602_ ;
wire \mylsu/_0603_ ;
wire \mylsu/_0604_ ;
wire \mylsu/_0605_ ;
wire \mylsu/_0606_ ;
wire \mylsu/_0607_ ;
wire \mylsu/_0608_ ;
wire \mylsu/_0609_ ;
wire \mylsu/_0610_ ;
wire \mylsu/_0611_ ;
wire \mylsu/_0612_ ;
wire \mylsu/_0613_ ;
wire \mylsu/_0614_ ;
wire \mylsu/_0615_ ;
wire \mylsu/_0616_ ;
wire \mylsu/_0617_ ;
wire \mylsu/_0618_ ;
wire \mylsu/_0619_ ;
wire \mylsu/_0620_ ;
wire \mylsu/_0621_ ;
wire \mylsu/_0622_ ;
wire \mylsu/_0623_ ;
wire \mylsu/_0624_ ;
wire \mylsu/_0625_ ;
wire \mylsu/_0626_ ;
wire \mylsu/_0627_ ;
wire \mylsu/_0628_ ;
wire \mylsu/_0629_ ;
wire \mylsu/_0630_ ;
wire \mylsu/_0631_ ;
wire \mylsu/_0632_ ;
wire \mylsu/_0633_ ;
wire \mylsu/_0634_ ;
wire \mylsu/_0635_ ;
wire \mylsu/_0636_ ;
wire \mylsu/_0637_ ;
wire \mylsu/_0638_ ;
wire \mylsu/_0639_ ;
wire \mylsu/_0640_ ;
wire \mylsu/_0641_ ;
wire \mylsu/_0642_ ;
wire \mylsu/_0643_ ;
wire \mylsu/_0644_ ;
wire \mylsu/_0645_ ;
wire \mylsu/_0646_ ;
wire \mylsu/_0647_ ;
wire \mylsu/_0648_ ;
wire \mylsu/_0649_ ;
wire \mylsu/_0650_ ;
wire \mylsu/_0651_ ;
wire \mylsu/_0652_ ;
wire \mylsu/_0653_ ;
wire \mylsu/_0654_ ;
wire \mylsu/_0655_ ;
wire \mylsu/_0656_ ;
wire \mylsu/_0657_ ;
wire \mylsu/_0658_ ;
wire \mylsu/_0659_ ;
wire \mylsu/_0660_ ;
wire \mylsu/_0661_ ;
wire \mylsu/_0662_ ;
wire \mylsu/_0663_ ;
wire \mylsu/_0664_ ;
wire \mylsu/_0665_ ;
wire \mylsu/_0666_ ;
wire \mylsu/_0667_ ;
wire \mylsu/_0668_ ;
wire \mylsu/_0669_ ;
wire \mylsu/_0670_ ;
wire \mylsu/_0671_ ;
wire \mylsu/_0672_ ;
wire \mylsu/_0673_ ;
wire \mylsu/_0674_ ;
wire \mylsu/_0675_ ;
wire \mylsu/_0676_ ;
wire \mylsu/_0677_ ;
wire \mylsu/_0678_ ;
wire \mylsu/_0679_ ;
wire \mylsu/_0680_ ;
wire \mylsu/_0681_ ;
wire \mylsu/_0682_ ;
wire \mylsu/_0683_ ;
wire \mylsu/_0684_ ;
wire \mylsu/_0685_ ;
wire \mylsu/_0686_ ;
wire \mylsu/_0687_ ;
wire \mylsu/_0688_ ;
wire \mylsu/_0689_ ;
wire \mylsu/_0690_ ;
wire \mylsu/_0691_ ;
wire \mylsu/_0692_ ;
wire \mylsu/_0693_ ;
wire \mylsu/_0694_ ;
wire \mylsu/_0695_ ;
wire \mylsu/_0696_ ;
wire \mylsu/_0697_ ;
wire \mylsu/_0698_ ;
wire \mylsu/_0699_ ;
wire \mylsu/_0700_ ;
wire \mylsu/_0701_ ;
wire \mylsu/_0702_ ;
wire \mylsu/_0703_ ;
wire \mylsu/_0704_ ;
wire \mylsu/_0705_ ;
wire \mylsu/_0706_ ;
wire \mylsu/_0707_ ;
wire \mylsu/_0708_ ;
wire \mylsu/_0709_ ;
wire \mylsu/_0710_ ;
wire \mylsu/_0711_ ;
wire \mylsu/_0712_ ;
wire \mylsu/_0713_ ;
wire \mylsu/_0714_ ;
wire \mylsu/_0715_ ;
wire \mylsu/_0716_ ;
wire \mylsu/_0717_ ;
wire \mylsu/_0718_ ;
wire \mylsu/_0719_ ;
wire \mylsu/_0720_ ;
wire \mylsu/_0721_ ;
wire \mylsu/_0722_ ;
wire \mylsu/_0723_ ;
wire \mylsu/_0724_ ;
wire \mylsu/_0725_ ;
wire \mylsu/_0726_ ;
wire \mylsu/_0727_ ;
wire \mylsu/_0728_ ;
wire \mylsu/_0729_ ;
wire \mylsu/_0730_ ;
wire \mylsu/_0731_ ;
wire \mylsu/_0732_ ;
wire \mylsu/_0733_ ;
wire \mylsu/_0734_ ;
wire \mylsu/_0735_ ;
wire \mylsu/_0736_ ;
wire \mylsu/_0737_ ;
wire \mylsu/_0738_ ;
wire \mylsu/_0739_ ;
wire \mylsu/_0740_ ;
wire \mylsu/_0741_ ;
wire \mylsu/_0742_ ;
wire \mylsu/_0743_ ;
wire \mylsu/_0744_ ;
wire \mylsu/_0745_ ;
wire \mylsu/_0746_ ;
wire \mylsu/_0747_ ;
wire \mylsu/_0748_ ;
wire \mylsu/_0749_ ;
wire \mylsu/_0750_ ;
wire \mylsu/_0751_ ;
wire \mylsu/_0752_ ;
wire \mylsu/_0753_ ;
wire \mylsu/_0754_ ;
wire \mylsu/_0755_ ;
wire \mylsu/_0756_ ;
wire \mylsu/_0757_ ;
wire \mylsu/_0758_ ;
wire \mylsu/_0759_ ;
wire \mylsu/_0760_ ;
wire \mylsu/_0761_ ;
wire \mylsu/_0762_ ;
wire \mylsu/_0763_ ;
wire \mylsu/_0764_ ;
wire \mylsu/_0765_ ;
wire \mylsu/_0766_ ;
wire \mylsu/_0767_ ;
wire \mylsu/_0768_ ;
wire \mylsu/_0769_ ;
wire \mylsu/_0770_ ;
wire \mylsu/_0771_ ;
wire \mylsu/_0772_ ;
wire \mylsu/_0773_ ;
wire \mylsu/_0774_ ;
wire \mylsu/_0775_ ;
wire \mylsu/_0776_ ;
wire \mylsu/_0777_ ;
wire \mylsu/_0778_ ;
wire \mylsu/_0779_ ;
wire \mylsu/_0780_ ;
wire \mylsu/_0781_ ;
wire \mylsu/_0782_ ;
wire \mylsu/_0783_ ;
wire \mylsu/_0784_ ;
wire \mylsu/_0785_ ;
wire \mylsu/_0786_ ;
wire \mylsu/_0787_ ;
wire \mylsu/_0788_ ;
wire \mylsu/_0789_ ;
wire \mylsu/_0790_ ;
wire \mylsu/_0791_ ;
wire \mylsu/_0792_ ;
wire \mylsu/_0793_ ;
wire \mylsu/_0794_ ;
wire \mylsu/_0795_ ;
wire \mylsu/_0796_ ;
wire \mylsu/_0797_ ;
wire \mylsu/_0798_ ;
wire \mylsu/_0799_ ;
wire \mylsu/_0800_ ;
wire \mylsu/_0801_ ;
wire \mylsu/_0802_ ;
wire \mylsu/_0803_ ;
wire \mylsu/_0804_ ;
wire \mylsu/_0805_ ;
wire \mylsu/_0806_ ;
wire \mylsu/_0807_ ;
wire \mylsu/_0808_ ;
wire \mylsu/_0809_ ;
wire \mylsu/_0810_ ;
wire \mylsu/_0811_ ;
wire \mylsu/_0812_ ;
wire \mylsu/_0813_ ;
wire \mylsu/_0814_ ;
wire \mylsu/_0815_ ;
wire \mylsu/_0816_ ;
wire \mylsu/_0817_ ;
wire \mylsu/_0818_ ;
wire \mylsu/_0819_ ;
wire \mylsu/_0820_ ;
wire \mylsu/_0821_ ;
wire \mylsu/_0822_ ;
wire \mylsu/_0823_ ;
wire \mylsu/_0824_ ;
wire \mylsu/_0825_ ;
wire \mylsu/_0826_ ;
wire \mylsu/_0827_ ;
wire \mylsu/_0828_ ;
wire \mylsu/_0829_ ;
wire \mylsu/_0830_ ;
wire \mylsu/_0831_ ;
wire \mylsu/_0832_ ;
wire \mylsu/_0833_ ;
wire \mylsu/_0834_ ;
wire \mylsu/_0835_ ;
wire \mylsu/_0836_ ;
wire \mylsu/_0837_ ;
wire \mylsu/_0838_ ;
wire \mylsu/_0839_ ;
wire \mylsu/_0840_ ;
wire \mylsu/_0841_ ;
wire \mylsu/_0842_ ;
wire \mylsu/_0843_ ;
wire \mylsu/_0844_ ;
wire \mylsu/_0845_ ;
wire \mylsu/_0846_ ;
wire \mylsu/_0847_ ;
wire \mylsu/_0848_ ;
wire \mylsu/_0849_ ;
wire \mylsu/_0850_ ;
wire \mylsu/_0851_ ;
wire \mylsu/_0852_ ;
wire \mylsu/_0853_ ;
wire \mylsu/_0854_ ;
wire \mylsu/_0855_ ;
wire \mylsu/_0856_ ;
wire \mylsu/_0857_ ;
wire \mylsu/_0858_ ;
wire \mylsu/_0859_ ;
wire \mylsu/_0860_ ;
wire \mylsu/_0861_ ;
wire \mylsu/_0862_ ;
wire \mylsu/_0863_ ;
wire \mylsu/_0864_ ;
wire \mylsu/_0865_ ;
wire \mylsu/_0866_ ;
wire \mylsu/_0867_ ;
wire \mylsu/_0868_ ;
wire \mylsu/_0869_ ;
wire \mylsu/_0870_ ;
wire \mylsu/_0871_ ;
wire \mylsu/_0872_ ;
wire \mylsu/_0873_ ;
wire \mylsu/_0874_ ;
wire \mylsu/_0875_ ;
wire \mylsu/_0876_ ;
wire \mylsu/_0877_ ;
wire \mylsu/_0878_ ;
wire \mylsu/_0879_ ;
wire \mylsu/_0880_ ;
wire \mylsu/_0881_ ;
wire \mylsu/_0882_ ;
wire \mylsu/_0883_ ;
wire \mylsu/_0884_ ;
wire \mylsu/_0885_ ;
wire \mylsu/_0886_ ;
wire \mylsu/_0887_ ;
wire \mylsu/_0888_ ;
wire \mylsu/_0889_ ;
wire \mylsu/_0890_ ;
wire \mylsu/_0891_ ;
wire \mylsu/_0892_ ;
wire \mylsu/_0893_ ;
wire \mylsu/_0894_ ;
wire \mylsu/_0895_ ;
wire \mylsu/_0896_ ;
wire \mylsu/_0897_ ;
wire \mylsu/_0898_ ;
wire \mylsu/_0899_ ;
wire \mylsu/_0900_ ;
wire \mylsu/_0901_ ;
wire \mylsu/_0902_ ;
wire \mylsu/_0903_ ;
wire \mylsu/_0904_ ;
wire \mylsu/_0905_ ;
wire \mylsu/_0906_ ;
wire \mylsu/_0907_ ;
wire \mylsu/_0908_ ;
wire \mylsu/_0909_ ;
wire \mylsu/_0910_ ;
wire \mylsu/_0911_ ;
wire \mylsu/_0912_ ;
wire \mylsu/_0913_ ;
wire \mylsu/_0914_ ;
wire \mylsu/_0915_ ;
wire \mylsu/_0916_ ;
wire \mylsu/_0917_ ;
wire \mylsu/_0918_ ;
wire \mylsu/_0919_ ;
wire \mylsu/_0920_ ;
wire \mylsu/_0921_ ;
wire \mylsu/_0922_ ;
wire \mylsu/_0923_ ;
wire \mylsu/_0924_ ;
wire \mylsu/_0925_ ;
wire \mylsu/_0926_ ;
wire \mylsu/_0927_ ;
wire \mylsu/_0928_ ;
wire \mylsu/_0929_ ;
wire \mylsu/_0930_ ;
wire \mylsu/_0931_ ;
wire \mylsu/_0932_ ;
wire \mylsu/_0933_ ;
wire \mylsu/_0934_ ;
wire \mylsu/_0935_ ;
wire \mylsu/_0936_ ;
wire \mylsu/_0937_ ;
wire \mylsu/_0938_ ;
wire \mylsu/_0939_ ;
wire \mylsu/_0940_ ;
wire \mylsu/_0941_ ;
wire \mylsu/_0942_ ;
wire \mylsu/_0943_ ;
wire \mylsu/_0944_ ;
wire \mylsu/_0945_ ;
wire \mylsu/_0946_ ;
wire \mylsu/_0947_ ;
wire \mylsu/_0948_ ;
wire \mylsu/_0949_ ;
wire \mylsu/_0950_ ;
wire \mylsu/_0951_ ;
wire \mylsu/_0952_ ;
wire \mylsu/_0953_ ;
wire \mylsu/_0954_ ;
wire \mylsu/_0955_ ;
wire \mylsu/_0956_ ;
wire \mylsu/_0957_ ;
wire \mylsu/_0958_ ;
wire \mylsu/_0959_ ;
wire \mylsu/_0960_ ;
wire \mylsu/_0961_ ;
wire \mylsu/_0962_ ;
wire \mylsu/_0963_ ;
wire \mylsu/_0964_ ;
wire \mylsu/_0965_ ;
wire \mylsu/_0966_ ;
wire \mylsu/_0967_ ;
wire \mylsu/_0968_ ;
wire \mylsu/_0969_ ;
wire \mylsu/_0970_ ;
wire \mylsu/_0971_ ;
wire \mylsu/_0972_ ;
wire \mylsu/_0973_ ;
wire \mylsu/_0974_ ;
wire \mylsu/_0975_ ;
wire \mylsu/_0976_ ;
wire \mylsu/_0977_ ;
wire \mylsu/_0978_ ;
wire \mylsu/_0979_ ;
wire \mylsu/_0980_ ;
wire \mylsu/_0981_ ;
wire \mylsu/_0982_ ;
wire \mylsu/_0983_ ;
wire \mylsu/_0984_ ;
wire \mylsu/_0985_ ;
wire \mylsu/_0986_ ;
wire \mylsu/_0987_ ;
wire \mylsu/_0988_ ;
wire \mylsu/_0989_ ;
wire \mylsu/_0990_ ;
wire \mylsu/_0991_ ;
wire \mylsu/_0992_ ;
wire \mylsu/_0993_ ;
wire \mylsu/_0994_ ;
wire \mylsu/_0995_ ;
wire \mylsu/_0996_ ;
wire \mylsu/_0997_ ;
wire \mylsu/_0998_ ;
wire \mylsu/_0999_ ;
wire \mylsu/_1000_ ;
wire \mylsu/_1001_ ;
wire \mylsu/_1002_ ;
wire \mylsu/_1003_ ;
wire \mylsu/_1004_ ;
wire \mylsu/_1005_ ;
wire \mylsu/_1006_ ;
wire \mylsu/_1007_ ;
wire \mylsu/_1008_ ;
wire \mylsu/_1009_ ;
wire \mylsu/_1010_ ;
wire \mylsu/_1011_ ;
wire \mylsu/_1012_ ;
wire \mylsu/_1013_ ;
wire \mylsu/_1014_ ;
wire \mylsu/_1015_ ;
wire \mylsu/_1016_ ;
wire \mylsu/_1017_ ;
wire \mylsu/_1018_ ;
wire \mylsu/_1019_ ;
wire \mylsu/_1020_ ;
wire \mylsu/_1021_ ;
wire \mylsu/_1022_ ;
wire \mylsu/_1023_ ;
wire \mylsu/_1024_ ;
wire \mylsu/_1025_ ;
wire \mylsu/_1026_ ;
wire \mylsu/_1027_ ;
wire \mylsu/_1028_ ;
wire \mylsu/_1029_ ;
wire \mylsu/_1030_ ;
wire \mylsu/_1031_ ;
wire \mylsu/_1032_ ;
wire \mylsu/_1033_ ;
wire \mylsu/_1034_ ;
wire \mylsu/_1035_ ;
wire \mylsu/_1036_ ;
wire \mylsu/_1037_ ;
wire \mylsu/_1038_ ;
wire \mylsu/_1039_ ;
wire \mylsu/_1040_ ;
wire \mylsu/_1041_ ;
wire \mylsu/_1042_ ;
wire \mylsu/_1043_ ;
wire \mylsu/_1044_ ;
wire \mylsu/_1045_ ;
wire \mylsu/_1046_ ;
wire \mylsu/_1047_ ;
wire \mylsu/_1048_ ;
wire \mylsu/_1049_ ;
wire \mylsu/_1050_ ;
wire \mylsu/_1051_ ;
wire \mylsu/_1052_ ;
wire \mylsu/_1053_ ;
wire \mylsu/_1054_ ;
wire \mylsu/_1055_ ;
wire \mylsu/_1056_ ;
wire \mylsu/_1057_ ;
wire \mylsu/_1058_ ;
wire \mylsu/_1059_ ;
wire \mylsu/_1060_ ;
wire \mylsu/_1061_ ;
wire \mylsu/_1062_ ;
wire \mylsu/_1063_ ;
wire \mylsu/_1064_ ;
wire \mylsu/_1065_ ;
wire \mylsu/_1066_ ;
wire \mylsu/_1067_ ;
wire \mylsu/_1068_ ;
wire \mylsu/_1069_ ;
wire \mylsu/_1070_ ;
wire \mylsu/_1071_ ;
wire \mylsu/_1072_ ;
wire \mylsu/_1073_ ;
wire \mylsu/_1074_ ;
wire \mylsu/_1075_ ;
wire \mylsu/_1076_ ;
wire \mylsu/_1077_ ;
wire \mylsu/_1078_ ;
wire \mylsu/_1079_ ;
wire \mylsu/_1080_ ;
wire \mylsu/_1081_ ;
wire \mylsu/_1082_ ;
wire \mylsu/_1083_ ;
wire \mylsu/_1084_ ;
wire \mylsu/_1085_ ;
wire \mylsu/_1086_ ;
wire \mylsu/_1087_ ;
wire \mylsu/_1088_ ;
wire \mylsu/_1089_ ;
wire \mylsu/_1090_ ;
wire \mylsu/_1091_ ;
wire \mylsu/_1092_ ;
wire \mylsu/_1093_ ;
wire \mylsu/_1094_ ;
wire \mylsu/_1095_ ;
wire \mylsu/_1096_ ;
wire \mylsu/_1097_ ;
wire \mylsu/_1098_ ;
wire \mylsu/_1099_ ;
wire \mylsu/_1100_ ;
wire \mylsu/_1101_ ;
wire \mylsu/_1102_ ;
wire \mylsu/_1103_ ;
wire \mylsu/_1104_ ;
wire \mylsu/_1105_ ;
wire \mylsu/_1106_ ;
wire \mylsu/_1107_ ;
wire \mylsu/_1108_ ;
wire \mylsu/_1109_ ;
wire \mylsu/_1110_ ;
wire \mylsu/_1111_ ;
wire \mylsu/_1112_ ;
wire \mylsu/_1113_ ;
wire \mylsu/_1114_ ;
wire \mylsu/_1115_ ;
wire \mylsu/_1116_ ;
wire \mylsu/_1117_ ;
wire \mylsu/_1118_ ;
wire \mylsu/_1119_ ;
wire \mylsu/_1120_ ;
wire \mylsu/_1121_ ;
wire \mylsu/_1122_ ;
wire \mylsu/_1123_ ;
wire \mylsu/_1124_ ;
wire \mylsu/_1125_ ;
wire \mylsu/_1126_ ;
wire \mylsu/_1127_ ;
wire \mylsu/_1128_ ;
wire \mylsu/_1129_ ;
wire \mylsu/_1130_ ;
wire \mylsu/_1131_ ;
wire \mylsu/_1132_ ;
wire \mylsu/_1133_ ;
wire \mylsu/_1134_ ;
wire \mylsu/_1135_ ;
wire \mylsu/_1136_ ;
wire \mylsu/_1137_ ;
wire \mylsu/_1138_ ;
wire \mylsu/_1139_ ;
wire \mylsu/_1140_ ;
wire \mylsu/_1141_ ;
wire \mylsu/_1142_ ;
wire \mylsu/_1143_ ;
wire \mylsu/_1144_ ;
wire \mylsu/_1145_ ;
wire \mylsu/_1146_ ;
wire \mylsu/_1147_ ;
wire \mylsu/_1148_ ;
wire \mylsu/_1149_ ;
wire \mylsu/_1150_ ;
wire \mylsu/_1151_ ;
wire \mylsu/_1152_ ;
wire \mylsu/_1153_ ;
wire \mylsu/_1154_ ;
wire \mylsu/_1155_ ;
wire \mylsu/_1156_ ;
wire \mylsu/_1157_ ;
wire \mylsu/_1158_ ;
wire \mylsu/_1159_ ;
wire \mylsu/_1160_ ;
wire \mylsu/_1161_ ;
wire \mylsu/_1162_ ;
wire \mylsu/_1163_ ;
wire \mylsu/_1164_ ;
wire \mylsu/_1165_ ;
wire \mylsu/_1166_ ;
wire \mylsu/_1167_ ;
wire \mylsu/_1168_ ;
wire \mylsu/_1169_ ;
wire \mylsu/_1170_ ;
wire \mylsu/_1171_ ;
wire \mylsu/_1172_ ;
wire \mylsu/_1173_ ;
wire \mylsu/_1174_ ;
wire \mylsu/_1175_ ;
wire \mylsu/_1176_ ;
wire \mylsu/_1177_ ;
wire \mylsu/_1178_ ;
wire \mylsu/_1179_ ;
wire \mylsu/_1180_ ;
wire \mylsu/_1181_ ;
wire \mylsu/_1182_ ;
wire \mylsu/_1183_ ;
wire \mylsu/_1184_ ;
wire \mylsu/_1185_ ;
wire \mylsu/_1186_ ;
wire \mylsu/_1187_ ;
wire \mylsu/_1188_ ;
wire \mylsu/_1189_ ;
wire \mylsu/_1190_ ;
wire \mylsu/_1191_ ;
wire \mylsu/_1192_ ;
wire \mylsu/_1193_ ;
wire \mylsu/_1194_ ;
wire \mylsu/_1195_ ;
wire \mylsu/_1196_ ;
wire \mylsu/_1197_ ;
wire \mylsu/_1198_ ;
wire \mylsu/_1199_ ;
wire \mylsu/_1200_ ;
wire \mylsu/_1201_ ;
wire \mylsu/_1202_ ;
wire \mylsu/_1203_ ;
wire \mylsu/_1204_ ;
wire \mylsu/_1205_ ;
wire \mylsu/_1206_ ;
wire \mylsu/_1207_ ;
wire \mylsu/_1208_ ;
wire \mylsu/_1209_ ;
wire \mylsu/_1210_ ;
wire \mylsu/_1211_ ;
wire \mylsu/_1212_ ;
wire \mylsu/_1213_ ;
wire \mylsu/_1214_ ;
wire \mylsu/_1215_ ;
wire \mylsu/_1216_ ;
wire \mylsu/_1217_ ;
wire \mylsu/_1218_ ;
wire \mylsu/_1219_ ;
wire \mylsu/_1220_ ;
wire \mylsu/_1221_ ;
wire \mylsu/_1222_ ;
wire \mylsu/_1223_ ;
wire \mylsu/_1224_ ;
wire \mylsu/_1225_ ;
wire \mylsu/_1226_ ;
wire \mylsu/_1227_ ;
wire \mylsu/_1228_ ;
wire \mylsu/_1229_ ;
wire \mylsu/_1230_ ;
wire \mylsu/_1231_ ;
wire \mylsu/_1232_ ;
wire \mylsu/_1233_ ;
wire \mylsu/_1234_ ;
wire \mylsu/_1235_ ;
wire \mylsu/_1236_ ;
wire \mylsu/_1237_ ;
wire \mylsu/_1238_ ;
wire \mylsu/_1239_ ;
wire \mylsu/_1240_ ;
wire \mylsu/_1241_ ;
wire \mylsu/_1242_ ;
wire \mylsu/_1243_ ;
wire \mylsu/_1244_ ;
wire \mylsu/_1245_ ;
wire \mylsu/_1246_ ;
wire \mylsu/_1247_ ;
wire \mylsu/_1248_ ;
wire \mylsu/_1249_ ;
wire \mylsu/_1250_ ;
wire \mylsu/_1251_ ;
wire \mylsu/_1252_ ;
wire \mylsu/_1253_ ;
wire \mylsu/_1254_ ;
wire \mylsu/_1255_ ;
wire \mylsu/_1256_ ;
wire \mylsu/_1257_ ;
wire \mylsu/_1258_ ;
wire \mylsu/_1259_ ;
wire \mylsu/_1260_ ;
wire \mylsu/_1261_ ;
wire \mylsu/_1262_ ;
wire \mylsu/_1263_ ;
wire \mylsu/_1264_ ;
wire \mylsu/_1265_ ;
wire \mylsu/_1266_ ;
wire \mylsu/_1267_ ;
wire \mylsu/_1268_ ;
wire \mylsu/_1269_ ;
wire \mylsu/_1270_ ;
wire \mylsu/_1271_ ;
wire \mylsu/_1272_ ;
wire \mylsu/_1273_ ;
wire \mylsu/_1274_ ;
wire \mylsu/_1275_ ;
wire \mylsu/_1276_ ;
wire \mylsu/_1277_ ;
wire \mylsu/_1278_ ;
wire \mylsu/_1279_ ;
wire \mylsu/_1280_ ;
wire \mylsu/_1281_ ;
wire \mylsu/_1282_ ;
wire \mylsu/_1283_ ;
wire \mylsu/_1284_ ;
wire \mylsu/_1285_ ;
wire \mylsu/_1286_ ;
wire \mylsu/_1287_ ;
wire \mylsu/_1288_ ;
wire \mylsu/_1289_ ;
wire \mylsu/_1290_ ;
wire \mylsu/_1291_ ;
wire \mylsu/_1292_ ;
wire \mylsu/_1293_ ;
wire \mylsu/_1294_ ;
wire \mylsu/_1295_ ;
wire \mylsu/_1296_ ;
wire \mylsu/_1297_ ;
wire \mylsu/_1298_ ;
wire \mylsu/_1299_ ;
wire \mylsu/_1300_ ;
wire \mylsu/_1301_ ;
wire \mylsu/_1302_ ;
wire \mylsu/_1303_ ;
wire \mylsu/_1304_ ;
wire \mylsu/_1305_ ;
wire \mylsu/_1306_ ;
wire \mylsu/_1307_ ;
wire \mylsu/_1308_ ;
wire \mylsu/_1309_ ;
wire \mylsu/_1310_ ;
wire \mylsu/_1311_ ;
wire \mylsu/_1312_ ;
wire \mylsu/_1313_ ;
wire \mylsu/_1314_ ;
wire \mylsu/_1315_ ;
wire \mylsu/_1316_ ;
wire \mylsu/_1317_ ;
wire \mylsu/_1318_ ;
wire \mylsu/_1319_ ;
wire \mylsu/_1320_ ;
wire \mylsu/_1321_ ;
wire \mylsu/_1322_ ;
wire \mylsu/_1323_ ;
wire \mylsu/_1324_ ;
wire \mylsu/_1325_ ;
wire \mylsu/_1326_ ;
wire \mylsu/_1327_ ;
wire \mylsu/_1328_ ;
wire \mylsu/_1329_ ;
wire \mylsu/_1330_ ;
wire \mylsu/_1331_ ;
wire \mylsu/_1332_ ;
wire \mylsu/_1333_ ;
wire \mylsu/_1334_ ;
wire \mylsu/_1335_ ;
wire \mylsu/_1336_ ;
wire \mylsu/_1337_ ;
wire \mylsu/_1338_ ;
wire \mylsu/_1339_ ;
wire \mylsu/_1340_ ;
wire \mylsu/_1341_ ;
wire \mylsu/_1342_ ;
wire \mylsu/_1343_ ;
wire \mylsu/_1344_ ;
wire \mylsu/_1345_ ;
wire \mylsu/_1346_ ;
wire \mylsu/_1347_ ;
wire \mylsu/_1348_ ;
wire \mylsu/_1349_ ;
wire \mylsu/_1350_ ;
wire \mylsu/_1351_ ;
wire \mylsu/_1352_ ;
wire \mylsu/_1353_ ;
wire \mylsu/_1354_ ;
wire \mylsu/_1355_ ;
wire \mylsu/_1356_ ;
wire \mylsu/_1357_ ;
wire \mylsu/_1358_ ;
wire \mylsu/_1359_ ;
wire \mylsu/_1360_ ;
wire \mylsu/_1361_ ;
wire \mylsu/_1362_ ;
wire \mylsu/_1363_ ;
wire \mylsu/_1364_ ;
wire \mylsu/_1365_ ;
wire \myminixbar/_0000_ ;
wire \myminixbar/_0001_ ;
wire \myminixbar/_0002_ ;
wire \myminixbar/_0003_ ;
wire \myminixbar/_0004_ ;
wire \myminixbar/_0005_ ;
wire \myminixbar/_0006_ ;
wire \myminixbar/_0007_ ;
wire \myminixbar/_0008_ ;
wire \myminixbar/_0009_ ;
wire \myminixbar/_0010_ ;
wire \myminixbar/_0011_ ;
wire \myminixbar/_0012_ ;
wire \myminixbar/_0013_ ;
wire \myminixbar/_0014_ ;
wire \myminixbar/_0015_ ;
wire \myminixbar/_0016_ ;
wire \myminixbar/_0017_ ;
wire \myminixbar/_0018_ ;
wire \myminixbar/_0019_ ;
wire \myminixbar/_0020_ ;
wire \myminixbar/_0021_ ;
wire \myminixbar/_0022_ ;
wire \myminixbar/_0023_ ;
wire \myminixbar/_0024_ ;
wire \myminixbar/_0025_ ;
wire \myminixbar/_0026_ ;
wire \myminixbar/_0027_ ;
wire \myminixbar/_0028_ ;
wire \myminixbar/_0029_ ;
wire \myminixbar/_0030_ ;
wire \myminixbar/_0031_ ;
wire \myminixbar/_0032_ ;
wire \myminixbar/_0033_ ;
wire \myminixbar/_0034_ ;
wire \myminixbar/_0035_ ;
wire \myminixbar/_0036_ ;
wire \myminixbar/_0037_ ;
wire \myminixbar/_0038_ ;
wire \myminixbar/_0039_ ;
wire \myminixbar/_0040_ ;
wire \myminixbar/_0041_ ;
wire \myminixbar/_0042_ ;
wire \myminixbar/_0043_ ;
wire \myminixbar/_0044_ ;
wire \myminixbar/_0045_ ;
wire \myminixbar/_0046_ ;
wire \myminixbar/_0047_ ;
wire \myminixbar/_0048_ ;
wire \myminixbar/_0049_ ;
wire \myminixbar/_0050_ ;
wire \myminixbar/_0051_ ;
wire \myminixbar/_0052_ ;
wire \myminixbar/_0053_ ;
wire \myminixbar/_0054_ ;
wire \myminixbar/_0055_ ;
wire \myminixbar/_0056_ ;
wire \myminixbar/_0057_ ;
wire \myminixbar/_0058_ ;
wire \myminixbar/_0059_ ;
wire \myminixbar/_0060_ ;
wire \myminixbar/_0061_ ;
wire \myminixbar/_0062_ ;
wire \myminixbar/_0063_ ;
wire \myminixbar/_0064_ ;
wire \myminixbar/_0065_ ;
wire \myminixbar/_0066_ ;
wire \myminixbar/_0067_ ;
wire \myminixbar/_0068_ ;
wire \myminixbar/_0069_ ;
wire \myminixbar/_0070_ ;
wire \myminixbar/_0071_ ;
wire \myminixbar/_0072_ ;
wire \myminixbar/_0073_ ;
wire \myminixbar/_0074_ ;
wire \myminixbar/_0075_ ;
wire \myminixbar/_0076_ ;
wire \myminixbar/_0077_ ;
wire \myminixbar/_0078_ ;
wire \myminixbar/_0079_ ;
wire \myminixbar/_0080_ ;
wire \myminixbar/_0081_ ;
wire \myminixbar/_0082_ ;
wire \myminixbar/_0083_ ;
wire \myminixbar/_0084_ ;
wire \myminixbar/_0085_ ;
wire \myminixbar/_0086_ ;
wire \myminixbar/_0087_ ;
wire \myminixbar/_0088_ ;
wire \myminixbar/_0089_ ;
wire \myminixbar/_0090_ ;
wire \myminixbar/_0091_ ;
wire \myminixbar/_0092_ ;
wire \myminixbar/_0093_ ;
wire \myminixbar/_0094_ ;
wire \myminixbar/_0095_ ;
wire \myminixbar/_0096_ ;
wire \myminixbar/_0097_ ;
wire \myminixbar/_0098_ ;
wire \myminixbar/_0099_ ;
wire \myminixbar/_0100_ ;
wire \myminixbar/_0101_ ;
wire \myminixbar/_0102_ ;
wire \myminixbar/_0103_ ;
wire \myminixbar/_0104_ ;
wire \myminixbar/_0105_ ;
wire \myminixbar/_0106_ ;
wire \myminixbar/_0107_ ;
wire \myminixbar/_0108_ ;
wire \myminixbar/_0109_ ;
wire \myminixbar/_0110_ ;
wire \myminixbar/_0111_ ;
wire \myminixbar/_0112_ ;
wire \myminixbar/_0113_ ;
wire \myminixbar/_0114_ ;
wire \myminixbar/_0115_ ;
wire \myminixbar/_0116_ ;
wire \myminixbar/_0117_ ;
wire \myminixbar/_0118_ ;
wire \myminixbar/_0119_ ;
wire \myminixbar/_0120_ ;
wire \myminixbar/_0121_ ;
wire \myminixbar/_0122_ ;
wire \myminixbar/_0123_ ;
wire \myminixbar/_0124_ ;
wire \myminixbar/_0125_ ;
wire \myminixbar/_0126_ ;
wire \myminixbar/_0127_ ;
wire \myminixbar/_0128_ ;
wire \myminixbar/_0129_ ;
wire \myminixbar/_0130_ ;
wire \myminixbar/_0131_ ;
wire \myminixbar/_0132_ ;
wire \myminixbar/_0133_ ;
wire \myminixbar/_0134_ ;
wire \myminixbar/_0135_ ;
wire \myminixbar/_0136_ ;
wire \myminixbar/_0137_ ;
wire \myminixbar/_0138_ ;
wire \myminixbar/_0139_ ;
wire \myminixbar/_0140_ ;
wire \myminixbar/_0141_ ;
wire \myminixbar/_0142_ ;
wire \myminixbar/_0143_ ;
wire \myminixbar/_0144_ ;
wire \myminixbar/_0145_ ;
wire \myminixbar/_0146_ ;
wire \myminixbar/_0147_ ;
wire \myminixbar/_0148_ ;
wire \myminixbar/_0149_ ;
wire \myminixbar/_0150_ ;
wire \myminixbar/_0151_ ;
wire \myminixbar/_0152_ ;
wire \myminixbar/_0153_ ;
wire \myminixbar/_0154_ ;
wire \myminixbar/_0155_ ;
wire \myminixbar/_0156_ ;
wire \myminixbar/_0157_ ;
wire \myminixbar/_0158_ ;
wire \myminixbar/_0159_ ;
wire \myminixbar/_0160_ ;
wire \myminixbar/_0161_ ;
wire \myminixbar/_0162_ ;
wire \myminixbar/_0163_ ;
wire \myminixbar/_0164_ ;
wire \myminixbar/_0165_ ;
wire \myminixbar/_0166_ ;
wire \myminixbar/_0167_ ;
wire \myminixbar/_0168_ ;
wire \myminixbar/_0169_ ;
wire \myminixbar/_0170_ ;
wire \myminixbar/_0171_ ;
wire \myminixbar/_0172_ ;
wire \myminixbar/_0173_ ;
wire \myminixbar/_0174_ ;
wire \myminixbar/_0175_ ;
wire \myminixbar/_0176_ ;
wire \myminixbar/_0177_ ;
wire \myminixbar/_0178_ ;
wire \myminixbar/_0179_ ;
wire \myminixbar/_0180_ ;
wire \myminixbar/_0181_ ;
wire \myminixbar/_0182_ ;
wire \myminixbar/_0183_ ;
wire \myminixbar/_0184_ ;
wire \myminixbar/_0185_ ;
wire \myminixbar/_0186_ ;
wire \myminixbar/_0187_ ;
wire \myminixbar/_0188_ ;
wire \myminixbar/_0189_ ;
wire \myminixbar/_0190_ ;
wire \myminixbar/_0191_ ;
wire \myminixbar/_0192_ ;
wire \myminixbar/_0193_ ;
wire \myminixbar/_0194_ ;
wire \myminixbar/_0195_ ;
wire \myminixbar/_0196_ ;
wire \myminixbar/_0197_ ;
wire \myminixbar/_0198_ ;
wire \myminixbar/_0199_ ;
wire \myminixbar/_0200_ ;
wire \myminixbar/_0201_ ;
wire \myminixbar/_0202_ ;
wire \myminixbar/_0203_ ;
wire \myminixbar/_0204_ ;
wire \myminixbar/_0205_ ;
wire \myminixbar/_0206_ ;
wire \myminixbar/_0207_ ;
wire \myminixbar/_0208_ ;
wire \myminixbar/_0209_ ;
wire \myminixbar/_0210_ ;
wire \myminixbar/_0211_ ;
wire \myminixbar/_0212_ ;
wire \myminixbar/_0213_ ;
wire \myminixbar/_0214_ ;
wire \myminixbar/_0215_ ;
wire \myminixbar/_0216_ ;
wire \myminixbar/_0217_ ;
wire \myminixbar/_0218_ ;
wire \myminixbar/_0219_ ;
wire \myminixbar/_0220_ ;
wire \myminixbar/_0221_ ;
wire \myminixbar/_0222_ ;
wire \myminixbar/_0223_ ;
wire \myminixbar/_0224_ ;
wire \myminixbar/_0225_ ;
wire \myminixbar/_0226_ ;
wire \myminixbar/_0227_ ;
wire \myminixbar/_0228_ ;
wire \myminixbar/_0229_ ;
wire \myminixbar/_0230_ ;
wire \myminixbar/_0231_ ;
wire \myminixbar/_0232_ ;
wire \myminixbar/_0233_ ;
wire \myminixbar/_0234_ ;
wire \myminixbar/_0235_ ;
wire \myminixbar/_0236_ ;
wire \myminixbar/_0237_ ;
wire \myminixbar/_0238_ ;
wire \myminixbar/_0239_ ;
wire \myminixbar/_0240_ ;
wire \myminixbar/_0241_ ;
wire \myminixbar/_0242_ ;
wire \myminixbar/_0243_ ;
wire \myminixbar/_0244_ ;
wire \myminixbar/_0245_ ;
wire \myminixbar/_0246_ ;
wire \myminixbar/_0247_ ;
wire \myminixbar/_0248_ ;
wire \myminixbar/_0249_ ;
wire \myminixbar/_0250_ ;
wire \myminixbar/_0251_ ;
wire \myminixbar/_0252_ ;
wire \myminixbar/_0253_ ;
wire \myminixbar/_0254_ ;
wire \myminixbar/_0255_ ;
wire \myminixbar/_0256_ ;
wire \myminixbar/_0257_ ;
wire \myminixbar/_0258_ ;
wire \myminixbar/_0259_ ;
wire \myminixbar/_0260_ ;
wire \myminixbar/_0261_ ;
wire \myminixbar/_0262_ ;
wire \myminixbar/_0263_ ;
wire \myminixbar/_0264_ ;
wire \myminixbar/_0265_ ;
wire \myminixbar/_0266_ ;
wire \myminixbar/_0267_ ;
wire \myminixbar/_0268_ ;
wire \myminixbar/_0269_ ;
wire \myminixbar/_0270_ ;
wire \myminixbar/_0271_ ;
wire \myminixbar/_0272_ ;
wire \myminixbar/_0273_ ;
wire \myminixbar/_0274_ ;
wire \myminixbar/_0275_ ;
wire \myminixbar/_0276_ ;
wire \myminixbar/_0277_ ;
wire \myminixbar/_0278_ ;
wire \myminixbar/_0279_ ;
wire \myminixbar/_0280_ ;
wire \myminixbar/_0281_ ;
wire \myminixbar/_0282_ ;
wire \myminixbar/_0283_ ;
wire \myminixbar/_0284_ ;
wire \myminixbar/_0285_ ;
wire \myminixbar/_0286_ ;
wire \myminixbar/_0287_ ;
wire \myminixbar/_0288_ ;
wire \myminixbar/_0289_ ;
wire \myminixbar/_0290_ ;
wire \myminixbar/_0291_ ;
wire \myminixbar/_0292_ ;
wire \myminixbar/_0293_ ;
wire \myminixbar/_0294_ ;
wire \myminixbar/_0295_ ;
wire \myminixbar/_0296_ ;
wire \myminixbar/_0297_ ;
wire \myminixbar/_0298_ ;
wire \myminixbar/_0299_ ;
wire \myminixbar/_0300_ ;
wire \myminixbar/_0301_ ;
wire \myminixbar/_0302_ ;
wire \myminixbar/_0303_ ;
wire \myminixbar/_0304_ ;
wire \myminixbar/_0305_ ;
wire \myminixbar/_0306_ ;
wire \myminixbar/_0307_ ;
wire \myminixbar/_0308_ ;
wire \myminixbar/_0309_ ;
wire \myminixbar/_0310_ ;
wire \myminixbar/_0311_ ;
wire \myminixbar/_0312_ ;
wire \myminixbar/_0313_ ;
wire \myminixbar/_0314_ ;
wire \myminixbar/_0315_ ;
wire \myminixbar/_0316_ ;
wire \myminixbar/_0317_ ;
wire \myminixbar/_0318_ ;
wire \myminixbar/_0319_ ;
wire \myminixbar/_0320_ ;
wire \myminixbar/_0321_ ;
wire \myminixbar/_0322_ ;
wire \myminixbar/_0323_ ;
wire \myminixbar/_0324_ ;
wire \myminixbar/_0325_ ;
wire \myminixbar/_0326_ ;
wire \myminixbar/_0327_ ;
wire \myminixbar/_0328_ ;
wire \myminixbar/_0329_ ;
wire \myminixbar/_0330_ ;
wire \myminixbar/_0331_ ;
wire \myminixbar/_0332_ ;
wire \myminixbar/_0333_ ;
wire \myminixbar/_0334_ ;
wire \myminixbar/_0335_ ;
wire \myminixbar/_0336_ ;
wire \myminixbar/_0337_ ;
wire \myminixbar/_0338_ ;
wire \myminixbar/_0339_ ;
wire \myminixbar/_0340_ ;
wire \myminixbar/_0341_ ;
wire \myminixbar/_0342_ ;
wire \myminixbar/_0343_ ;
wire \myminixbar/_0344_ ;
wire \myminixbar/_0345_ ;
wire \myminixbar/_0346_ ;
wire \myminixbar/_0347_ ;
wire \myminixbar/_0348_ ;
wire \myminixbar/_0349_ ;
wire \myminixbar/_0350_ ;
wire \myminixbar/_0351_ ;
wire \myminixbar/_0352_ ;
wire \myminixbar/_0353_ ;
wire \myminixbar/_0354_ ;
wire \myminixbar/_0355_ ;
wire \myminixbar/_0356_ ;
wire \myminixbar/_0357_ ;
wire \myminixbar/_0358_ ;
wire \myminixbar/_0359_ ;
wire \myminixbar/_0360_ ;
wire \myminixbar/_0361_ ;
wire \myminixbar/_0362_ ;
wire \myminixbar/_0363_ ;
wire \myminixbar/_0364_ ;
wire \myminixbar/_0365_ ;
wire \myminixbar/_0366_ ;
wire \myminixbar/_0367_ ;
wire \myminixbar/_0368_ ;
wire \myminixbar/_0369_ ;
wire \myminixbar/_0370_ ;
wire \myminixbar/_0371_ ;
wire \myminixbar/_0372_ ;
wire \myminixbar/_0373_ ;
wire \myminixbar/_0374_ ;
wire \myminixbar/_0375_ ;
wire \myminixbar/_0376_ ;
wire \myminixbar/_0377_ ;
wire \myminixbar/_0378_ ;
wire \myminixbar/_0379_ ;
wire \myminixbar/_0380_ ;
wire \myminixbar/_0381_ ;
wire \myminixbar/_0382_ ;
wire \myminixbar/_0383_ ;
wire \myminixbar/_0384_ ;
wire \myminixbar/_0385_ ;
wire \myminixbar/_0386_ ;
wire \myminixbar/_0387_ ;
wire \myminixbar/_0388_ ;
wire \myminixbar/_0389_ ;
wire \myminixbar/_0390_ ;
wire \myminixbar/_0391_ ;
wire \myminixbar/_0392_ ;
wire \myminixbar/_0393_ ;
wire \myminixbar/_0394_ ;
wire \myminixbar/_0395_ ;
wire \myminixbar/_0396_ ;
wire \myminixbar/_0397_ ;
wire \myminixbar/_0398_ ;
wire \myminixbar/_0399_ ;
wire \myminixbar/_0400_ ;
wire \myminixbar/_0401_ ;
wire \myminixbar/_0402_ ;
wire \myminixbar/_0403_ ;
wire \myminixbar/_0404_ ;
wire \myminixbar/_0405_ ;
wire \myminixbar/_0406_ ;
wire \myminixbar/_0407_ ;
wire \myminixbar/_0408_ ;
wire \myminixbar/_0409_ ;
wire \myminixbar/_0410_ ;
wire \myminixbar/_0411_ ;
wire \myminixbar/_0412_ ;
wire \myminixbar/_0413_ ;
wire \myminixbar/_0414_ ;
wire \myminixbar/_0415_ ;
wire \myminixbar/_0416_ ;
wire \myminixbar/_0417_ ;
wire \myminixbar/_0418_ ;
wire \myminixbar/_0419_ ;
wire \myminixbar/_0420_ ;
wire \myminixbar/_0421_ ;
wire \myminixbar/_0422_ ;
wire \myminixbar/_0423_ ;
wire \myminixbar/_0424_ ;
wire \myminixbar/_0425_ ;
wire \myminixbar/_0426_ ;
wire \myminixbar/_0427_ ;
wire \myminixbar/_0428_ ;
wire \myminixbar/_0429_ ;
wire \myminixbar/_0430_ ;
wire \myminixbar/_0431_ ;
wire \myminixbar/_0432_ ;
wire \myminixbar/_0433_ ;
wire \myminixbar/_0434_ ;
wire \myminixbar/_0435_ ;
wire \myminixbar/_0436_ ;
wire \myminixbar/_0437_ ;
wire \myminixbar/_0438_ ;
wire \myminixbar/_0439_ ;
wire \myminixbar/_0440_ ;
wire \myminixbar/_0441_ ;
wire \myminixbar/_0442_ ;
wire \myminixbar/_0443_ ;
wire \myminixbar/_0444_ ;
wire \myminixbar/_0445_ ;
wire \myminixbar/_0446_ ;
wire \myminixbar/_0447_ ;
wire \myminixbar/_0448_ ;
wire \myminixbar/_0449_ ;
wire \myminixbar/_0450_ ;
wire \myminixbar/_0451_ ;
wire \myminixbar/_0452_ ;
wire \myminixbar/_0453_ ;
wire \myminixbar/_0454_ ;
wire \myminixbar/_0455_ ;
wire \myminixbar/_0456_ ;
wire \myminixbar/_0457_ ;
wire \myminixbar/_0458_ ;
wire \myminixbar/_0459_ ;
wire \myminixbar/_0460_ ;
wire \myminixbar/_0461_ ;
wire \myminixbar/_0462_ ;
wire \myminixbar/_0463_ ;
wire \myminixbar/_0464_ ;
wire \myminixbar/_0465_ ;
wire \myminixbar/_0466_ ;
wire \myminixbar/_0467_ ;
wire \myminixbar/_0468_ ;
wire \myminixbar/_0469_ ;
wire \myminixbar/_0470_ ;
wire \myminixbar/_0471_ ;
wire \myminixbar/_0472_ ;
wire \myminixbar/_0473_ ;
wire \myminixbar/_0474_ ;
wire \myminixbar/_0475_ ;
wire \myminixbar/_0476_ ;
wire \myminixbar/_0477_ ;
wire \myminixbar/_0478_ ;
wire \myminixbar/_0479_ ;
wire \myminixbar/_0480_ ;
wire \myminixbar/_0481_ ;
wire \myminixbar/_0482_ ;
wire \myminixbar/_0483_ ;
wire \myminixbar/_0484_ ;
wire \myminixbar/_0485_ ;
wire \myminixbar/_0486_ ;
wire \myminixbar/_0487_ ;
wire \myminixbar/_0488_ ;
wire \myminixbar/_0489_ ;
wire \myminixbar/_0490_ ;
wire \myminixbar/_0491_ ;
wire \myminixbar/_0492_ ;
wire \myminixbar/_0493_ ;
wire \myminixbar/_0494_ ;
wire \myminixbar/_0495_ ;
wire \myminixbar/_0496_ ;
wire \myminixbar/_0497_ ;
wire \myminixbar/_0498_ ;
wire \myminixbar/_0499_ ;
wire \myminixbar/_0500_ ;
wire \myminixbar/_0501_ ;
wire \myminixbar/_0502_ ;
wire \myminixbar/_0503_ ;
wire \myminixbar/_0504_ ;
wire \myminixbar/_0505_ ;
wire \myminixbar/_0506_ ;
wire \myminixbar/_0507_ ;
wire \myreg/_0000_ ;
wire \myreg/_0001_ ;
wire \myreg/_0002_ ;
wire \myreg/_0003_ ;
wire \myreg/_0004_ ;
wire \myreg/_0005_ ;
wire \myreg/_0006_ ;
wire \myreg/_0007_ ;
wire \myreg/_0008_ ;
wire \myreg/_0009_ ;
wire \myreg/_0010_ ;
wire \myreg/_0011_ ;
wire \myreg/_0012_ ;
wire \myreg/_0013_ ;
wire \myreg/_0014_ ;
wire \myreg/_0015_ ;
wire \myreg/_0016_ ;
wire \myreg/_0017_ ;
wire \myreg/_0018_ ;
wire \myreg/_0019_ ;
wire \myreg/_0020_ ;
wire \myreg/_0021_ ;
wire \myreg/_0022_ ;
wire \myreg/_0023_ ;
wire \myreg/_0024_ ;
wire \myreg/_0025_ ;
wire \myreg/_0026_ ;
wire \myreg/_0027_ ;
wire \myreg/_0028_ ;
wire \myreg/_0029_ ;
wire \myreg/_0030_ ;
wire \myreg/_0031_ ;
wire \myreg/_0032_ ;
wire \myreg/_0033_ ;
wire \myreg/_0034_ ;
wire \myreg/_0035_ ;
wire \myreg/_0036_ ;
wire \myreg/_0037_ ;
wire \myreg/_0038_ ;
wire \myreg/_0039_ ;
wire \myreg/_0040_ ;
wire \myreg/_0041_ ;
wire \myreg/_0042_ ;
wire \myreg/_0043_ ;
wire \myreg/_0044_ ;
wire \myreg/_0045_ ;
wire \myreg/_0046_ ;
wire \myreg/_0047_ ;
wire \myreg/_0048_ ;
wire \myreg/_0049_ ;
wire \myreg/_0050_ ;
wire \myreg/_0051_ ;
wire \myreg/_0052_ ;
wire \myreg/_0053_ ;
wire \myreg/_0054_ ;
wire \myreg/_0055_ ;
wire \myreg/_0056_ ;
wire \myreg/_0057_ ;
wire \myreg/_0058_ ;
wire \myreg/_0059_ ;
wire \myreg/_0060_ ;
wire \myreg/_0061_ ;
wire \myreg/_0062_ ;
wire \myreg/_0063_ ;
wire \myreg/_0064_ ;
wire \myreg/_0065_ ;
wire \myreg/_0066_ ;
wire \myreg/_0067_ ;
wire \myreg/_0068_ ;
wire \myreg/_0069_ ;
wire \myreg/_0070_ ;
wire \myreg/_0071_ ;
wire \myreg/_0072_ ;
wire \myreg/_0073_ ;
wire \myreg/_0074_ ;
wire \myreg/_0075_ ;
wire \myreg/_0076_ ;
wire \myreg/_0077_ ;
wire \myreg/_0078_ ;
wire \myreg/_0079_ ;
wire \myreg/_0080_ ;
wire \myreg/_0081_ ;
wire \myreg/_0082_ ;
wire \myreg/_0083_ ;
wire \myreg/_0084_ ;
wire \myreg/_0085_ ;
wire \myreg/_0086_ ;
wire \myreg/_0087_ ;
wire \myreg/_0088_ ;
wire \myreg/_0089_ ;
wire \myreg/_0090_ ;
wire \myreg/_0091_ ;
wire \myreg/_0092_ ;
wire \myreg/_0093_ ;
wire \myreg/_0094_ ;
wire \myreg/_0095_ ;
wire \myreg/_0096_ ;
wire \myreg/_0097_ ;
wire \myreg/_0098_ ;
wire \myreg/_0099_ ;
wire \myreg/_0100_ ;
wire \myreg/_0101_ ;
wire \myreg/_0102_ ;
wire \myreg/_0103_ ;
wire \myreg/_0104_ ;
wire \myreg/_0105_ ;
wire \myreg/_0106_ ;
wire \myreg/_0107_ ;
wire \myreg/_0108_ ;
wire \myreg/_0109_ ;
wire \myreg/_0110_ ;
wire \myreg/_0111_ ;
wire \myreg/_0112_ ;
wire \myreg/_0113_ ;
wire \myreg/_0114_ ;
wire \myreg/_0115_ ;
wire \myreg/_0116_ ;
wire \myreg/_0117_ ;
wire \myreg/_0118_ ;
wire \myreg/_0119_ ;
wire \myreg/_0120_ ;
wire \myreg/_0121_ ;
wire \myreg/_0122_ ;
wire \myreg/_0123_ ;
wire \myreg/_0124_ ;
wire \myreg/_0125_ ;
wire \myreg/_0126_ ;
wire \myreg/_0127_ ;
wire \myreg/_0128_ ;
wire \myreg/_0129_ ;
wire \myreg/_0130_ ;
wire \myreg/_0131_ ;
wire \myreg/_0132_ ;
wire \myreg/_0133_ ;
wire \myreg/_0134_ ;
wire \myreg/_0135_ ;
wire \myreg/_0136_ ;
wire \myreg/_0137_ ;
wire \myreg/_0138_ ;
wire \myreg/_0139_ ;
wire \myreg/_0140_ ;
wire \myreg/_0141_ ;
wire \myreg/_0142_ ;
wire \myreg/_0143_ ;
wire \myreg/_0144_ ;
wire \myreg/_0145_ ;
wire \myreg/_0146_ ;
wire \myreg/_0147_ ;
wire \myreg/_0148_ ;
wire \myreg/_0149_ ;
wire \myreg/_0150_ ;
wire \myreg/_0151_ ;
wire \myreg/_0152_ ;
wire \myreg/_0153_ ;
wire \myreg/_0154_ ;
wire \myreg/_0155_ ;
wire \myreg/_0156_ ;
wire \myreg/_0157_ ;
wire \myreg/_0158_ ;
wire \myreg/_0159_ ;
wire \myreg/_0160_ ;
wire \myreg/_0161_ ;
wire \myreg/_0162_ ;
wire \myreg/_0163_ ;
wire \myreg/_0164_ ;
wire \myreg/_0165_ ;
wire \myreg/_0166_ ;
wire \myreg/_0167_ ;
wire \myreg/_0168_ ;
wire \myreg/_0169_ ;
wire \myreg/_0170_ ;
wire \myreg/_0171_ ;
wire \myreg/_0172_ ;
wire \myreg/_0173_ ;
wire \myreg/_0174_ ;
wire \myreg/_0175_ ;
wire \myreg/_0176_ ;
wire \myreg/_0177_ ;
wire \myreg/_0178_ ;
wire \myreg/_0179_ ;
wire \myreg/_0180_ ;
wire \myreg/_0181_ ;
wire \myreg/_0182_ ;
wire \myreg/_0183_ ;
wire \myreg/_0184_ ;
wire \myreg/_0185_ ;
wire \myreg/_0186_ ;
wire \myreg/_0187_ ;
wire \myreg/_0188_ ;
wire \myreg/_0189_ ;
wire \myreg/_0190_ ;
wire \myreg/_0191_ ;
wire \myreg/_0192_ ;
wire \myreg/_0193_ ;
wire \myreg/_0194_ ;
wire \myreg/_0195_ ;
wire \myreg/_0196_ ;
wire \myreg/_0197_ ;
wire \myreg/_0198_ ;
wire \myreg/_0199_ ;
wire \myreg/_0200_ ;
wire \myreg/_0201_ ;
wire \myreg/_0202_ ;
wire \myreg/_0203_ ;
wire \myreg/_0204_ ;
wire \myreg/_0205_ ;
wire \myreg/_0206_ ;
wire \myreg/_0207_ ;
wire \myreg/_0208_ ;
wire \myreg/_0209_ ;
wire \myreg/_0210_ ;
wire \myreg/_0211_ ;
wire \myreg/_0212_ ;
wire \myreg/_0213_ ;
wire \myreg/_0214_ ;
wire \myreg/_0215_ ;
wire \myreg/_0216_ ;
wire \myreg/_0217_ ;
wire \myreg/_0218_ ;
wire \myreg/_0219_ ;
wire \myreg/_0220_ ;
wire \myreg/_0221_ ;
wire \myreg/_0222_ ;
wire \myreg/_0223_ ;
wire \myreg/_0224_ ;
wire \myreg/_0225_ ;
wire \myreg/_0226_ ;
wire \myreg/_0227_ ;
wire \myreg/_0228_ ;
wire \myreg/_0229_ ;
wire \myreg/_0230_ ;
wire \myreg/_0231_ ;
wire \myreg/_0232_ ;
wire \myreg/_0233_ ;
wire \myreg/_0234_ ;
wire \myreg/_0235_ ;
wire \myreg/_0236_ ;
wire \myreg/_0237_ ;
wire \myreg/_0238_ ;
wire \myreg/_0239_ ;
wire \myreg/_0240_ ;
wire \myreg/_0241_ ;
wire \myreg/_0242_ ;
wire \myreg/_0243_ ;
wire \myreg/_0244_ ;
wire \myreg/_0245_ ;
wire \myreg/_0246_ ;
wire \myreg/_0247_ ;
wire \myreg/_0248_ ;
wire \myreg/_0249_ ;
wire \myreg/_0250_ ;
wire \myreg/_0251_ ;
wire \myreg/_0252_ ;
wire \myreg/_0253_ ;
wire \myreg/_0254_ ;
wire \myreg/_0255_ ;
wire \myreg/_0256_ ;
wire \myreg/_0257_ ;
wire \myreg/_0258_ ;
wire \myreg/_0259_ ;
wire \myreg/_0260_ ;
wire \myreg/_0261_ ;
wire \myreg/_0262_ ;
wire \myreg/_0263_ ;
wire \myreg/_0264_ ;
wire \myreg/_0265_ ;
wire \myreg/_0266_ ;
wire \myreg/_0267_ ;
wire \myreg/_0268_ ;
wire \myreg/_0269_ ;
wire \myreg/_0270_ ;
wire \myreg/_0271_ ;
wire \myreg/_0272_ ;
wire \myreg/_0273_ ;
wire \myreg/_0274_ ;
wire \myreg/_0275_ ;
wire \myreg/_0276_ ;
wire \myreg/_0277_ ;
wire \myreg/_0278_ ;
wire \myreg/_0279_ ;
wire \myreg/_0280_ ;
wire \myreg/_0281_ ;
wire \myreg/_0282_ ;
wire \myreg/_0283_ ;
wire \myreg/_0284_ ;
wire \myreg/_0285_ ;
wire \myreg/_0286_ ;
wire \myreg/_0287_ ;
wire \myreg/_0288_ ;
wire \myreg/_0289_ ;
wire \myreg/_0290_ ;
wire \myreg/_0291_ ;
wire \myreg/_0292_ ;
wire \myreg/_0293_ ;
wire \myreg/_0294_ ;
wire \myreg/_0295_ ;
wire \myreg/_0296_ ;
wire \myreg/_0297_ ;
wire \myreg/_0298_ ;
wire \myreg/_0299_ ;
wire \myreg/_0300_ ;
wire \myreg/_0301_ ;
wire \myreg/_0302_ ;
wire \myreg/_0303_ ;
wire \myreg/_0304_ ;
wire \myreg/_0305_ ;
wire \myreg/_0306_ ;
wire \myreg/_0307_ ;
wire \myreg/_0308_ ;
wire \myreg/_0309_ ;
wire \myreg/_0310_ ;
wire \myreg/_0311_ ;
wire \myreg/_0312_ ;
wire \myreg/_0313_ ;
wire \myreg/_0314_ ;
wire \myreg/_0315_ ;
wire \myreg/_0316_ ;
wire \myreg/_0317_ ;
wire \myreg/_0318_ ;
wire \myreg/_0319_ ;
wire \myreg/_0320_ ;
wire \myreg/_0321_ ;
wire \myreg/_0322_ ;
wire \myreg/_0323_ ;
wire \myreg/_0324_ ;
wire \myreg/_0325_ ;
wire \myreg/_0326_ ;
wire \myreg/_0327_ ;
wire \myreg/_0328_ ;
wire \myreg/_0329_ ;
wire \myreg/_0330_ ;
wire \myreg/_0331_ ;
wire \myreg/_0332_ ;
wire \myreg/_0333_ ;
wire \myreg/_0334_ ;
wire \myreg/_0335_ ;
wire \myreg/_0336_ ;
wire \myreg/_0337_ ;
wire \myreg/_0338_ ;
wire \myreg/_0339_ ;
wire \myreg/_0340_ ;
wire \myreg/_0341_ ;
wire \myreg/_0342_ ;
wire \myreg/_0343_ ;
wire \myreg/_0344_ ;
wire \myreg/_0345_ ;
wire \myreg/_0346_ ;
wire \myreg/_0347_ ;
wire \myreg/_0348_ ;
wire \myreg/_0349_ ;
wire \myreg/_0350_ ;
wire \myreg/_0351_ ;
wire \myreg/_0352_ ;
wire \myreg/_0353_ ;
wire \myreg/_0354_ ;
wire \myreg/_0355_ ;
wire \myreg/_0356_ ;
wire \myreg/_0357_ ;
wire \myreg/_0358_ ;
wire \myreg/_0359_ ;
wire \myreg/_0360_ ;
wire \myreg/_0361_ ;
wire \myreg/_0362_ ;
wire \myreg/_0363_ ;
wire \myreg/_0364_ ;
wire \myreg/_0365_ ;
wire \myreg/_0366_ ;
wire \myreg/_0367_ ;
wire \myreg/_0368_ ;
wire \myreg/_0369_ ;
wire \myreg/_0370_ ;
wire \myreg/_0371_ ;
wire \myreg/_0372_ ;
wire \myreg/_0373_ ;
wire \myreg/_0374_ ;
wire \myreg/_0375_ ;
wire \myreg/_0376_ ;
wire \myreg/_0377_ ;
wire \myreg/_0378_ ;
wire \myreg/_0379_ ;
wire \myreg/_0380_ ;
wire \myreg/_0381_ ;
wire \myreg/_0382_ ;
wire \myreg/_0383_ ;
wire \myreg/_0384_ ;
wire \myreg/_0385_ ;
wire \myreg/_0386_ ;
wire \myreg/_0387_ ;
wire \myreg/_0388_ ;
wire \myreg/_0389_ ;
wire \myreg/_0390_ ;
wire \myreg/_0391_ ;
wire \myreg/_0392_ ;
wire \myreg/_0393_ ;
wire \myreg/_0394_ ;
wire \myreg/_0395_ ;
wire \myreg/_0396_ ;
wire \myreg/_0397_ ;
wire \myreg/_0398_ ;
wire \myreg/_0399_ ;
wire \myreg/_0400_ ;
wire \myreg/_0401_ ;
wire \myreg/_0402_ ;
wire \myreg/_0403_ ;
wire \myreg/_0404_ ;
wire \myreg/_0405_ ;
wire \myreg/_0406_ ;
wire \myreg/_0407_ ;
wire \myreg/_0408_ ;
wire \myreg/_0409_ ;
wire \myreg/_0410_ ;
wire \myreg/_0411_ ;
wire \myreg/_0412_ ;
wire \myreg/_0413_ ;
wire \myreg/_0414_ ;
wire \myreg/_0415_ ;
wire \myreg/_0416_ ;
wire \myreg/_0417_ ;
wire \myreg/_0418_ ;
wire \myreg/_0419_ ;
wire \myreg/_0420_ ;
wire \myreg/_0421_ ;
wire \myreg/_0422_ ;
wire \myreg/_0423_ ;
wire \myreg/_0424_ ;
wire \myreg/_0425_ ;
wire \myreg/_0426_ ;
wire \myreg/_0427_ ;
wire \myreg/_0428_ ;
wire \myreg/_0429_ ;
wire \myreg/_0430_ ;
wire \myreg/_0431_ ;
wire \myreg/_0432_ ;
wire \myreg/_0433_ ;
wire \myreg/_0434_ ;
wire \myreg/_0435_ ;
wire \myreg/_0436_ ;
wire \myreg/_0437_ ;
wire \myreg/_0438_ ;
wire \myreg/_0439_ ;
wire \myreg/_0440_ ;
wire \myreg/_0441_ ;
wire \myreg/_0442_ ;
wire \myreg/_0443_ ;
wire \myreg/_0444_ ;
wire \myreg/_0445_ ;
wire \myreg/_0446_ ;
wire \myreg/_0447_ ;
wire \myreg/_0448_ ;
wire \myreg/_0449_ ;
wire \myreg/_0450_ ;
wire \myreg/_0451_ ;
wire \myreg/_0452_ ;
wire \myreg/_0453_ ;
wire \myreg/_0454_ ;
wire \myreg/_0455_ ;
wire \myreg/_0456_ ;
wire \myreg/_0457_ ;
wire \myreg/_0458_ ;
wire \myreg/_0459_ ;
wire \myreg/_0460_ ;
wire \myreg/_0461_ ;
wire \myreg/_0462_ ;
wire \myreg/_0463_ ;
wire \myreg/_0464_ ;
wire \myreg/_0465_ ;
wire \myreg/_0466_ ;
wire \myreg/_0467_ ;
wire \myreg/_0468_ ;
wire \myreg/_0469_ ;
wire \myreg/_0470_ ;
wire \myreg/_0471_ ;
wire \myreg/_0472_ ;
wire \myreg/_0473_ ;
wire \myreg/_0474_ ;
wire \myreg/_0475_ ;
wire \myreg/_0476_ ;
wire \myreg/_0477_ ;
wire \myreg/_0478_ ;
wire \myreg/_0479_ ;
wire \myreg/_0480_ ;
wire \myreg/_0481_ ;
wire \myreg/_0482_ ;
wire \myreg/_0483_ ;
wire \myreg/_0484_ ;
wire \myreg/_0485_ ;
wire \myreg/_0486_ ;
wire \myreg/_0487_ ;
wire \myreg/_0488_ ;
wire \myreg/_0489_ ;
wire \myreg/_0490_ ;
wire \myreg/_0491_ ;
wire \myreg/_0492_ ;
wire \myreg/_0493_ ;
wire \myreg/_0494_ ;
wire \myreg/_0495_ ;
wire \myreg/_0496_ ;
wire \myreg/_0497_ ;
wire \myreg/_0498_ ;
wire \myreg/_0499_ ;
wire \myreg/_0500_ ;
wire \myreg/_0501_ ;
wire \myreg/_0502_ ;
wire \myreg/_0503_ ;
wire \myreg/_0504_ ;
wire \myreg/_0505_ ;
wire \myreg/_0506_ ;
wire \myreg/_0507_ ;
wire \myreg/_0508_ ;
wire \myreg/_0509_ ;
wire \myreg/_0510_ ;
wire \myreg/_0511_ ;
wire \myreg/_0512_ ;
wire \myreg/_0513_ ;
wire \myreg/_0514_ ;
wire \myreg/_0515_ ;
wire \myreg/_0516_ ;
wire \myreg/_0517_ ;
wire \myreg/_0518_ ;
wire \myreg/_0519_ ;
wire \myreg/_0520_ ;
wire \myreg/_0521_ ;
wire \myreg/_0522_ ;
wire \myreg/_0523_ ;
wire \myreg/_0524_ ;
wire \myreg/_0525_ ;
wire \myreg/_0526_ ;
wire \myreg/_0527_ ;
wire \myreg/_0528_ ;
wire \myreg/_0529_ ;
wire \myreg/_0530_ ;
wire \myreg/_0531_ ;
wire \myreg/_0532_ ;
wire \myreg/_0533_ ;
wire \myreg/_0534_ ;
wire \myreg/_0535_ ;
wire \myreg/_0536_ ;
wire \myreg/_0537_ ;
wire \myreg/_0538_ ;
wire \myreg/_0539_ ;
wire \myreg/_0540_ ;
wire \myreg/_0541_ ;
wire \myreg/_0542_ ;
wire \myreg/_0543_ ;
wire \myreg/_0544_ ;
wire \myreg/_0545_ ;
wire \myreg/_0546_ ;
wire \myreg/_0547_ ;
wire \myreg/_0548_ ;
wire \myreg/_0549_ ;
wire \myreg/_0550_ ;
wire \myreg/_0551_ ;
wire \myreg/_0552_ ;
wire \myreg/_0553_ ;
wire \myreg/_0554_ ;
wire \myreg/_0555_ ;
wire \myreg/_0556_ ;
wire \myreg/_0557_ ;
wire \myreg/_0558_ ;
wire \myreg/_0559_ ;
wire \myreg/_0560_ ;
wire \myreg/_0561_ ;
wire \myreg/_0562_ ;
wire \myreg/_0563_ ;
wire \myreg/_0564_ ;
wire \myreg/_0565_ ;
wire \myreg/_0566_ ;
wire \myreg/_0567_ ;
wire \myreg/_0568_ ;
wire \myreg/_0569_ ;
wire \myreg/_0570_ ;
wire \myreg/_0571_ ;
wire \myreg/_0572_ ;
wire \myreg/_0573_ ;
wire \myreg/_0574_ ;
wire \myreg/_0575_ ;
wire \myreg/_0576_ ;
wire \myreg/_0577_ ;
wire \myreg/_0578_ ;
wire \myreg/_0579_ ;
wire \myreg/_0580_ ;
wire \myreg/_0581_ ;
wire \myreg/_0582_ ;
wire \myreg/_0583_ ;
wire \myreg/_0584_ ;
wire \myreg/_0585_ ;
wire \myreg/_0586_ ;
wire \myreg/_0587_ ;
wire \myreg/_0588_ ;
wire \myreg/_0589_ ;
wire \myreg/_0590_ ;
wire \myreg/_0591_ ;
wire \myreg/_0592_ ;
wire \myreg/_0593_ ;
wire \myreg/_0594_ ;
wire \myreg/_0595_ ;
wire \myreg/_0596_ ;
wire \myreg/_0597_ ;
wire \myreg/_0598_ ;
wire \myreg/_0599_ ;
wire \myreg/_0600_ ;
wire \myreg/_0601_ ;
wire \myreg/_0602_ ;
wire \myreg/_0603_ ;
wire \myreg/_0604_ ;
wire \myreg/_0605_ ;
wire \myreg/_0606_ ;
wire \myreg/_0607_ ;
wire \myreg/_0608_ ;
wire \myreg/_0609_ ;
wire \myreg/_0610_ ;
wire \myreg/_0611_ ;
wire \myreg/_0612_ ;
wire \myreg/_0613_ ;
wire \myreg/_0614_ ;
wire \myreg/_0615_ ;
wire \myreg/_0616_ ;
wire \myreg/_0617_ ;
wire \myreg/_0618_ ;
wire \myreg/_0619_ ;
wire \myreg/_0620_ ;
wire \myreg/_0621_ ;
wire \myreg/_0622_ ;
wire \myreg/_0623_ ;
wire \myreg/_0624_ ;
wire \myreg/_0625_ ;
wire \myreg/_0626_ ;
wire \myreg/_0627_ ;
wire \myreg/_0628_ ;
wire \myreg/_0629_ ;
wire \myreg/_0630_ ;
wire \myreg/_0631_ ;
wire \myreg/_0632_ ;
wire \myreg/_0633_ ;
wire \myreg/_0634_ ;
wire \myreg/_0635_ ;
wire \myreg/_0636_ ;
wire \myreg/_0637_ ;
wire \myreg/_0638_ ;
wire \myreg/_0639_ ;
wire \myreg/_0640_ ;
wire \myreg/_0641_ ;
wire \myreg/_0642_ ;
wire \myreg/_0643_ ;
wire \myreg/_0644_ ;
wire \myreg/_0645_ ;
wire \myreg/_0646_ ;
wire \myreg/_0647_ ;
wire \myreg/_0648_ ;
wire \myreg/_0649_ ;
wire \myreg/_0650_ ;
wire \myreg/_0651_ ;
wire \myreg/_0652_ ;
wire \myreg/_0653_ ;
wire \myreg/_0654_ ;
wire \myreg/_0655_ ;
wire \myreg/_0656_ ;
wire \myreg/_0657_ ;
wire \myreg/_0658_ ;
wire \myreg/_0659_ ;
wire \myreg/_0660_ ;
wire \myreg/_0661_ ;
wire \myreg/_0662_ ;
wire \myreg/_0663_ ;
wire \myreg/_0664_ ;
wire \myreg/_0665_ ;
wire \myreg/_0666_ ;
wire \myreg/_0667_ ;
wire \myreg/_0668_ ;
wire \myreg/_0669_ ;
wire \myreg/_0670_ ;
wire \myreg/_0671_ ;
wire \myreg/_0672_ ;
wire \myreg/_0673_ ;
wire \myreg/_0674_ ;
wire \myreg/_0675_ ;
wire \myreg/_0676_ ;
wire \myreg/_0677_ ;
wire \myreg/_0678_ ;
wire \myreg/_0679_ ;
wire \myreg/_0680_ ;
wire \myreg/_0681_ ;
wire \myreg/_0682_ ;
wire \myreg/_0683_ ;
wire \myreg/_0684_ ;
wire \myreg/_0685_ ;
wire \myreg/_0686_ ;
wire \myreg/_0687_ ;
wire \myreg/_0688_ ;
wire \myreg/_0689_ ;
wire \myreg/_0690_ ;
wire \myreg/_0691_ ;
wire \myreg/_0692_ ;
wire \myreg/_0693_ ;
wire \myreg/_0694_ ;
wire \myreg/_0695_ ;
wire \myreg/_0696_ ;
wire \myreg/_0697_ ;
wire \myreg/_0698_ ;
wire \myreg/_0699_ ;
wire \myreg/_0700_ ;
wire \myreg/_0701_ ;
wire \myreg/_0702_ ;
wire \myreg/_0703_ ;
wire \myreg/_0704_ ;
wire \myreg/_0705_ ;
wire \myreg/_0706_ ;
wire \myreg/_0707_ ;
wire \myreg/_0708_ ;
wire \myreg/_0709_ ;
wire \myreg/_0710_ ;
wire \myreg/_0711_ ;
wire \myreg/_0712_ ;
wire \myreg/_0713_ ;
wire \myreg/_0714_ ;
wire \myreg/_0715_ ;
wire \myreg/_0716_ ;
wire \myreg/_0717_ ;
wire \myreg/_0718_ ;
wire \myreg/_0719_ ;
wire \myreg/_0720_ ;
wire \myreg/_0721_ ;
wire \myreg/_0722_ ;
wire \myreg/_0723_ ;
wire \myreg/_0724_ ;
wire \myreg/_0725_ ;
wire \myreg/_0726_ ;
wire \myreg/_0727_ ;
wire \myreg/_0728_ ;
wire \myreg/_0729_ ;
wire \myreg/_0730_ ;
wire \myreg/_0731_ ;
wire \myreg/_0732_ ;
wire \myreg/_0733_ ;
wire \myreg/_0734_ ;
wire \myreg/_0735_ ;
wire \myreg/_0736_ ;
wire \myreg/_0737_ ;
wire \myreg/_0738_ ;
wire \myreg/_0739_ ;
wire \myreg/_0740_ ;
wire \myreg/_0741_ ;
wire \myreg/_0742_ ;
wire \myreg/_0743_ ;
wire \myreg/_0744_ ;
wire \myreg/_0745_ ;
wire \myreg/_0746_ ;
wire \myreg/_0747_ ;
wire \myreg/_0748_ ;
wire \myreg/_0749_ ;
wire \myreg/_0750_ ;
wire \myreg/_0751_ ;
wire \myreg/_0752_ ;
wire \myreg/_0753_ ;
wire \myreg/_0754_ ;
wire \myreg/_0755_ ;
wire \myreg/_0756_ ;
wire \myreg/_0757_ ;
wire \myreg/_0758_ ;
wire \myreg/_0759_ ;
wire \myreg/_0760_ ;
wire \myreg/_0761_ ;
wire \myreg/_0762_ ;
wire \myreg/_0763_ ;
wire \myreg/_0764_ ;
wire \myreg/_0765_ ;
wire \myreg/_0766_ ;
wire \myreg/_0767_ ;
wire \myreg/_0768_ ;
wire \myreg/_0769_ ;
wire \myreg/_0770_ ;
wire \myreg/_0771_ ;
wire \myreg/_0772_ ;
wire \myreg/_0773_ ;
wire \myreg/_0774_ ;
wire \myreg/_0775_ ;
wire \myreg/_0776_ ;
wire \myreg/_0777_ ;
wire \myreg/_0778_ ;
wire \myreg/_0779_ ;
wire \myreg/_0780_ ;
wire \myreg/_0781_ ;
wire \myreg/_0782_ ;
wire \myreg/_0783_ ;
wire \myreg/_0784_ ;
wire \myreg/_0785_ ;
wire \myreg/_0786_ ;
wire \myreg/_0787_ ;
wire \myreg/_0788_ ;
wire \myreg/_0789_ ;
wire \myreg/_0790_ ;
wire \myreg/_0791_ ;
wire \myreg/_0792_ ;
wire \myreg/_0793_ ;
wire \myreg/_0794_ ;
wire \myreg/_0795_ ;
wire \myreg/_0796_ ;
wire \myreg/_0797_ ;
wire \myreg/_0798_ ;
wire \myreg/_0799_ ;
wire \myreg/_0800_ ;
wire \myreg/_0801_ ;
wire \myreg/_0802_ ;
wire \myreg/_0803_ ;
wire \myreg/_0804_ ;
wire \myreg/_0805_ ;
wire \myreg/_0806_ ;
wire \myreg/_0807_ ;
wire \myreg/_0808_ ;
wire \myreg/_0809_ ;
wire \myreg/_0810_ ;
wire \myreg/_0811_ ;
wire \myreg/_0812_ ;
wire \myreg/_0813_ ;
wire \myreg/_0814_ ;
wire \myreg/_0815_ ;
wire \myreg/_0816_ ;
wire \myreg/_0817_ ;
wire \myreg/_0818_ ;
wire \myreg/_0819_ ;
wire \myreg/_0820_ ;
wire \myreg/_0821_ ;
wire \myreg/_0822_ ;
wire \myreg/_0823_ ;
wire \myreg/_0824_ ;
wire \myreg/_0825_ ;
wire \myreg/_0826_ ;
wire \myreg/_0827_ ;
wire \myreg/_0828_ ;
wire \myreg/_0829_ ;
wire \myreg/_0830_ ;
wire \myreg/_0831_ ;
wire \myreg/_0832_ ;
wire \myreg/_0833_ ;
wire \myreg/_0834_ ;
wire \myreg/_0835_ ;
wire \myreg/_0836_ ;
wire \myreg/_0837_ ;
wire \myreg/_0838_ ;
wire \myreg/_0839_ ;
wire \myreg/_0840_ ;
wire \myreg/_0841_ ;
wire \myreg/_0842_ ;
wire \myreg/_0843_ ;
wire \myreg/_0844_ ;
wire \myreg/_0845_ ;
wire \myreg/_0846_ ;
wire \myreg/_0847_ ;
wire \myreg/_0848_ ;
wire \myreg/_0849_ ;
wire \myreg/_0850_ ;
wire \myreg/_0851_ ;
wire \myreg/_0852_ ;
wire \myreg/_0853_ ;
wire \myreg/_0854_ ;
wire \myreg/_0855_ ;
wire \myreg/_0856_ ;
wire \myreg/_0857_ ;
wire \myreg/_0858_ ;
wire \myreg/_0859_ ;
wire \myreg/_0860_ ;
wire \myreg/_0861_ ;
wire \myreg/_0862_ ;
wire \myreg/_0863_ ;
wire \myreg/_0864_ ;
wire \myreg/_0865_ ;
wire \myreg/_0866_ ;
wire \myreg/_0867_ ;
wire \myreg/_0868_ ;
wire \myreg/_0869_ ;
wire \myreg/_0870_ ;
wire \myreg/_0871_ ;
wire \myreg/_0872_ ;
wire \myreg/_0873_ ;
wire \myreg/_0874_ ;
wire \myreg/_0875_ ;
wire \myreg/_0876_ ;
wire \myreg/_0877_ ;
wire \myreg/_0878_ ;
wire \myreg/_0879_ ;
wire \myreg/_0880_ ;
wire \myreg/_0881_ ;
wire \myreg/_0882_ ;
wire \myreg/_0883_ ;
wire \myreg/_0884_ ;
wire \myreg/_0885_ ;
wire \myreg/_0886_ ;
wire \myreg/_0887_ ;
wire \myreg/_0888_ ;
wire \myreg/_0889_ ;
wire \myreg/_0890_ ;
wire \myreg/_0891_ ;
wire \myreg/_0892_ ;
wire \myreg/_0893_ ;
wire \myreg/_0894_ ;
wire \myreg/_0895_ ;
wire \myreg/_0896_ ;
wire \myreg/_0897_ ;
wire \myreg/_0898_ ;
wire \myreg/_0899_ ;
wire \myreg/_0900_ ;
wire \myreg/_0901_ ;
wire \myreg/_0902_ ;
wire \myreg/_0903_ ;
wire \myreg/_0904_ ;
wire \myreg/_0905_ ;
wire \myreg/_0906_ ;
wire \myreg/_0907_ ;
wire \myreg/_0908_ ;
wire \myreg/_0909_ ;
wire \myreg/_0910_ ;
wire \myreg/_0911_ ;
wire \myreg/_0912_ ;
wire \myreg/_0913_ ;
wire \myreg/_0914_ ;
wire \myreg/_0915_ ;
wire \myreg/_0916_ ;
wire \myreg/_0917_ ;
wire \myreg/_0918_ ;
wire \myreg/_0919_ ;
wire \myreg/_0920_ ;
wire \myreg/_0921_ ;
wire \myreg/_0922_ ;
wire \myreg/_0923_ ;
wire \myreg/_0924_ ;
wire \myreg/_0925_ ;
wire \myreg/_0926_ ;
wire \myreg/_0927_ ;
wire \myreg/_0928_ ;
wire \myreg/_0929_ ;
wire \myreg/_0930_ ;
wire \myreg/_0931_ ;
wire \myreg/_0932_ ;
wire \myreg/_0933_ ;
wire \myreg/_0934_ ;
wire \myreg/_0935_ ;
wire \myreg/_0936_ ;
wire \myreg/_0937_ ;
wire \myreg/_0938_ ;
wire \myreg/_0939_ ;
wire \myreg/_0940_ ;
wire \myreg/_0941_ ;
wire \myreg/_0942_ ;
wire \myreg/_0943_ ;
wire \myreg/_0944_ ;
wire \myreg/_0945_ ;
wire \myreg/_0946_ ;
wire \myreg/_0947_ ;
wire \myreg/_0948_ ;
wire \myreg/_0949_ ;
wire \myreg/_0950_ ;
wire \myreg/_0951_ ;
wire \myreg/_0952_ ;
wire \myreg/_0953_ ;
wire \myreg/_0954_ ;
wire \myreg/_0955_ ;
wire \myreg/_0956_ ;
wire \myreg/_0957_ ;
wire \myreg/_0958_ ;
wire \myreg/_0959_ ;
wire \myreg/_0960_ ;
wire \myreg/_0961_ ;
wire \myreg/_0962_ ;
wire \myreg/_0963_ ;
wire \myreg/_0964_ ;
wire \myreg/_0965_ ;
wire \myreg/_0966_ ;
wire \myreg/_0967_ ;
wire \myreg/_0968_ ;
wire \myreg/_0969_ ;
wire \myreg/_0970_ ;
wire \myreg/_0971_ ;
wire \myreg/_0972_ ;
wire \myreg/_0973_ ;
wire \myreg/_0974_ ;
wire \myreg/_0975_ ;
wire \myreg/_0976_ ;
wire \myreg/_0977_ ;
wire \myreg/_0978_ ;
wire \myreg/_0979_ ;
wire \myreg/_0980_ ;
wire \myreg/_0981_ ;
wire \myreg/_0982_ ;
wire \myreg/_0983_ ;
wire \myreg/_0984_ ;
wire \myreg/_0985_ ;
wire \myreg/_0986_ ;
wire \myreg/_0987_ ;
wire \myreg/_0988_ ;
wire \myreg/_0989_ ;
wire \myreg/_0990_ ;
wire \myreg/_0991_ ;
wire \myreg/_0992_ ;
wire \myreg/_0993_ ;
wire \myreg/_0994_ ;
wire \myreg/_0995_ ;
wire \myreg/_0996_ ;
wire \myreg/_0997_ ;
wire \myreg/_0998_ ;
wire \myreg/_0999_ ;
wire \myreg/_1000_ ;
wire \myreg/_1001_ ;
wire \myreg/_1002_ ;
wire \myreg/_1003_ ;
wire \myreg/_1004_ ;
wire \myreg/_1005_ ;
wire \myreg/_1006_ ;
wire \myreg/_1007_ ;
wire \myreg/_1008_ ;
wire \myreg/_1009_ ;
wire \myreg/_1010_ ;
wire \myreg/_1011_ ;
wire \myreg/_1012_ ;
wire \myreg/_1013_ ;
wire \myreg/_1014_ ;
wire \myreg/_1015_ ;
wire \myreg/_1016_ ;
wire \myreg/_1017_ ;
wire \myreg/_1018_ ;
wire \myreg/_1019_ ;
wire \myreg/_1020_ ;
wire \myreg/_1021_ ;
wire \myreg/_1022_ ;
wire \myreg/_1023_ ;
wire \myreg/_1024_ ;
wire \myreg/_1025_ ;
wire \myreg/_1026_ ;
wire \myreg/_1027_ ;
wire \myreg/_1028_ ;
wire \myreg/_1029_ ;
wire \myreg/_1030_ ;
wire \myreg/_1031_ ;
wire \myreg/_1032_ ;
wire \myreg/_1033_ ;
wire \myreg/_1034_ ;
wire \myreg/_1035_ ;
wire \myreg/_1036_ ;
wire \myreg/_1037_ ;
wire \myreg/_1038_ ;
wire \myreg/_1039_ ;
wire \myreg/_1040_ ;
wire \myreg/_1041_ ;
wire \myreg/_1042_ ;
wire \myreg/_1043_ ;
wire \myreg/_1044_ ;
wire \myreg/_1045_ ;
wire \myreg/_1046_ ;
wire \myreg/_1047_ ;
wire \myreg/_1048_ ;
wire \myreg/_1049_ ;
wire \myreg/_1050_ ;
wire \myreg/_1051_ ;
wire \myreg/_1052_ ;
wire \myreg/_1053_ ;
wire \myreg/_1054_ ;
wire \myreg/_1055_ ;
wire \myreg/_1056_ ;
wire \myreg/_1057_ ;
wire \myreg/_1058_ ;
wire \myreg/_1059_ ;
wire \myreg/_1060_ ;
wire \myreg/_1061_ ;
wire \myreg/_1062_ ;
wire \myreg/_1063_ ;
wire \myreg/_1064_ ;
wire \myreg/_1065_ ;
wire \myreg/_1066_ ;
wire \myreg/_1067_ ;
wire \myreg/_1068_ ;
wire \myreg/_1069_ ;
wire \myreg/_1070_ ;
wire \myreg/_1071_ ;
wire \myreg/_1072_ ;
wire \myreg/_1073_ ;
wire \myreg/_1074_ ;
wire \myreg/_1075_ ;
wire \myreg/_1076_ ;
wire \myreg/_1077_ ;
wire \myreg/_1078_ ;
wire \myreg/_1079_ ;
wire \myreg/_1080_ ;
wire \myreg/_1081_ ;
wire \myreg/_1082_ ;
wire \myreg/_1083_ ;
wire \myreg/_1084_ ;
wire \myreg/_1085_ ;
wire \myreg/_1086_ ;
wire \myreg/_1087_ ;
wire \myreg/_1088_ ;
wire \myreg/_1089_ ;
wire \myreg/_1090_ ;
wire \myreg/_1091_ ;
wire \myreg/_1092_ ;
wire \myreg/_1093_ ;
wire \myreg/_1094_ ;
wire \myreg/_1095_ ;
wire \myreg/_1096_ ;
wire \myreg/_1097_ ;
wire \myreg/_1098_ ;
wire \myreg/_1099_ ;
wire \myreg/_1100_ ;
wire \myreg/_1101_ ;
wire \myreg/_1102_ ;
wire \myreg/_1103_ ;
wire \myreg/_1104_ ;
wire \myreg/_1105_ ;
wire \myreg/_1106_ ;
wire \myreg/_1107_ ;
wire \myreg/_1108_ ;
wire \myreg/_1109_ ;
wire \myreg/_1110_ ;
wire \myreg/_1111_ ;
wire \myreg/_1112_ ;
wire \myreg/_1113_ ;
wire \myreg/_1114_ ;
wire \myreg/_1115_ ;
wire \myreg/_1116_ ;
wire \myreg/_1117_ ;
wire \myreg/_1118_ ;
wire \myreg/_1119_ ;
wire \myreg/_1120_ ;
wire \myreg/_1121_ ;
wire \myreg/_1122_ ;
wire \myreg/_1123_ ;
wire \myreg/_1124_ ;
wire \myreg/_1125_ ;
wire \myreg/_1126_ ;
wire \myreg/_1127_ ;
wire \myreg/_1128_ ;
wire \myreg/_1129_ ;
wire \myreg/_1130_ ;
wire \myreg/_1131_ ;
wire \myreg/_1132_ ;
wire \myreg/_1133_ ;
wire \myreg/_1134_ ;
wire \myreg/_1135_ ;
wire \myreg/_1136_ ;
wire \myreg/_1137_ ;
wire \myreg/_1138_ ;
wire \myreg/_1139_ ;
wire \myreg/_1140_ ;
wire \myreg/_1141_ ;
wire \myreg/_1142_ ;
wire \myreg/_1143_ ;
wire \myreg/_1144_ ;
wire \myreg/_1145_ ;
wire \myreg/_1146_ ;
wire \myreg/_1147_ ;
wire \myreg/_1148_ ;
wire \myreg/_1149_ ;
wire \myreg/_1150_ ;
wire \myreg/_1151_ ;
wire \myreg/_1152_ ;
wire \myreg/_1153_ ;
wire \myreg/_1154_ ;
wire \myreg/_1155_ ;
wire \myreg/_1156_ ;
wire \myreg/_1157_ ;
wire \myreg/_1158_ ;
wire \myreg/_1159_ ;
wire \myreg/_1160_ ;
wire \myreg/_1161_ ;
wire \myreg/_1162_ ;
wire \myreg/_1163_ ;
wire \myreg/_1164_ ;
wire \myreg/_1165_ ;
wire \myreg/_1166_ ;
wire \myreg/_1167_ ;
wire \myreg/_1168_ ;
wire \myreg/_1169_ ;
wire \myreg/_1170_ ;
wire \myreg/_1171_ ;
wire \myreg/_1172_ ;
wire \myreg/_1173_ ;
wire \myreg/_1174_ ;
wire \myreg/_1175_ ;
wire \myreg/_1176_ ;
wire \myreg/_1177_ ;
wire \myreg/_1178_ ;
wire \myreg/_1179_ ;
wire \myreg/_1180_ ;
wire \myreg/_1181_ ;
wire \myreg/_1182_ ;
wire \myreg/_1183_ ;
wire \myreg/_1184_ ;
wire \myreg/_1185_ ;
wire \myreg/_1186_ ;
wire \myreg/_1187_ ;
wire \myreg/_1188_ ;
wire \myreg/_1189_ ;
wire \myreg/_1190_ ;
wire \myreg/_1191_ ;
wire \myreg/_1192_ ;
wire \myreg/_1193_ ;
wire \myreg/_1194_ ;
wire \myreg/_1195_ ;
wire \myreg/_1196_ ;
wire \myreg/_1197_ ;
wire \myreg/_1198_ ;
wire \myreg/_1199_ ;
wire \myreg/_1200_ ;
wire \myreg/_1201_ ;
wire \myreg/_1202_ ;
wire \myreg/_1203_ ;
wire \myreg/_1204_ ;
wire \myreg/_1205_ ;
wire \myreg/_1206_ ;
wire \myreg/_1207_ ;
wire \myreg/_1208_ ;
wire \myreg/_1209_ ;
wire \myreg/_1210_ ;
wire \myreg/_1211_ ;
wire \myreg/_1212_ ;
wire \myreg/_1213_ ;
wire \myreg/_1214_ ;
wire \myreg/_1215_ ;
wire \myreg/_1216_ ;
wire \myreg/_1217_ ;
wire \myreg/_1218_ ;
wire \myreg/_1219_ ;
wire \myreg/_1220_ ;
wire \myreg/_1221_ ;
wire \myreg/_1222_ ;
wire \myreg/_1223_ ;
wire \myreg/_1224_ ;
wire \myreg/_1225_ ;
wire \myreg/_1226_ ;
wire \myreg/_1227_ ;
wire \myreg/_1228_ ;
wire \myreg/_1229_ ;
wire \myreg/_1230_ ;
wire \myreg/_1231_ ;
wire \myreg/_1232_ ;
wire \myreg/_1233_ ;
wire \myreg/_1234_ ;
wire \myreg/_1235_ ;
wire \myreg/_1236_ ;
wire \myreg/_1237_ ;
wire \myreg/_1238_ ;
wire \myreg/_1239_ ;
wire \myreg/_1240_ ;
wire \myreg/_1241_ ;
wire \myreg/_1242_ ;
wire \myreg/_1243_ ;
wire \myreg/_1244_ ;
wire \myreg/_1245_ ;
wire \myreg/_1246_ ;
wire \myreg/_1247_ ;
wire \myreg/_1248_ ;
wire \myreg/_1249_ ;
wire \myreg/_1250_ ;
wire \myreg/_1251_ ;
wire \myreg/_1252_ ;
wire \myreg/_1253_ ;
wire \myreg/_1254_ ;
wire \myreg/_1255_ ;
wire \myreg/_1256_ ;
wire \myreg/_1257_ ;
wire \myreg/_1258_ ;
wire \myreg/_1259_ ;
wire \myreg/_1260_ ;
wire \myreg/_1261_ ;
wire \myreg/_1262_ ;
wire \myreg/_1263_ ;
wire \myreg/_1264_ ;
wire \myreg/_1265_ ;
wire \myreg/_1266_ ;
wire \myreg/_1267_ ;
wire \myreg/_1268_ ;
wire \myreg/_1269_ ;
wire \myreg/_1270_ ;
wire \myreg/_1271_ ;
wire \myreg/_1272_ ;
wire \myreg/_1273_ ;
wire \myreg/_1274_ ;
wire \myreg/_1275_ ;
wire \myreg/_1276_ ;
wire \myreg/_1277_ ;
wire \myreg/_1278_ ;
wire \myreg/_1279_ ;
wire \myreg/_1280_ ;
wire \myreg/_1281_ ;
wire \myreg/_1282_ ;
wire \myreg/_1283_ ;
wire \myreg/_1284_ ;
wire \myreg/_1285_ ;
wire \myreg/_1286_ ;
wire \myreg/_1287_ ;
wire \myreg/_1288_ ;
wire \myreg/_1289_ ;
wire \myreg/_1290_ ;
wire \myreg/_1291_ ;
wire \myreg/_1292_ ;
wire \myreg/_1293_ ;
wire \myreg/_1294_ ;
wire \myreg/_1295_ ;
wire \myreg/_1296_ ;
wire \myreg/_1297_ ;
wire \myreg/_1298_ ;
wire \myreg/_1299_ ;
wire \myreg/_1300_ ;
wire \myreg/_1301_ ;
wire \myreg/_1302_ ;
wire \myreg/_1303_ ;
wire \myreg/_1304_ ;
wire \myreg/_1305_ ;
wire \myreg/_1306_ ;
wire \myreg/_1307_ ;
wire \myreg/_1308_ ;
wire \myreg/_1309_ ;
wire \myreg/_1310_ ;
wire \myreg/_1311_ ;
wire \myreg/_1312_ ;
wire \myreg/_1313_ ;
wire \myreg/_1314_ ;
wire \myreg/_1315_ ;
wire \myreg/_1316_ ;
wire \myreg/_1317_ ;
wire \myreg/_1318_ ;
wire \myreg/_1319_ ;
wire \myreg/_1320_ ;
wire \myreg/_1321_ ;
wire \myreg/_1322_ ;
wire \myreg/_1323_ ;
wire \myreg/_1324_ ;
wire \myreg/_1325_ ;
wire \myreg/_1326_ ;
wire \myreg/_1327_ ;
wire \myreg/_1328_ ;
wire \myreg/_1329_ ;
wire \myreg/_1330_ ;
wire \myreg/_1331_ ;
wire \myreg/_1332_ ;
wire \myreg/_1333_ ;
wire \myreg/_1334_ ;
wire \myreg/_1335_ ;
wire \myreg/_1336_ ;
wire \myreg/_1337_ ;
wire \myreg/_1338_ ;
wire \myreg/_1339_ ;
wire \myreg/_1340_ ;
wire \myreg/_1341_ ;
wire \myreg/_1342_ ;
wire \myreg/_1343_ ;
wire \myreg/_1344_ ;
wire \myreg/_1345_ ;
wire \myreg/_1346_ ;
wire \myreg/_1347_ ;
wire \myreg/_1348_ ;
wire \myreg/_1349_ ;
wire \myreg/_1350_ ;
wire \myreg/_1351_ ;
wire \myreg/_1352_ ;
wire \myreg/_1353_ ;
wire \myreg/_1354_ ;
wire \myreg/_1355_ ;
wire \myreg/_1356_ ;
wire \myreg/_1357_ ;
wire \myreg/_1358_ ;
wire \myreg/_1359_ ;
wire \myreg/_1360_ ;
wire \myreg/_1361_ ;
wire \myreg/_1362_ ;
wire \myreg/_1363_ ;
wire \myreg/_1364_ ;
wire \myreg/_1365_ ;
wire \myreg/_1366_ ;
wire \myreg/_1367_ ;
wire \myreg/_1368_ ;
wire \myreg/_1369_ ;
wire \myreg/_1370_ ;
wire \myreg/_1371_ ;
wire \myreg/_1372_ ;
wire \myreg/_1373_ ;
wire \myreg/_1374_ ;
wire \myreg/_1375_ ;
wire \myreg/_1376_ ;
wire \myreg/_1377_ ;
wire \myreg/_1378_ ;
wire \myreg/_1379_ ;
wire \myreg/_1380_ ;
wire \myreg/_1381_ ;
wire \myreg/_1382_ ;
wire \myreg/_1383_ ;
wire \myreg/_1384_ ;
wire \myreg/_1385_ ;
wire \myreg/_1386_ ;
wire \myreg/_1387_ ;
wire \myreg/_1388_ ;
wire \myreg/_1389_ ;
wire \myreg/_1390_ ;
wire \myreg/_1391_ ;
wire \myreg/_1392_ ;
wire \myreg/_1393_ ;
wire \myreg/_1394_ ;
wire \myreg/_1395_ ;
wire \myreg/_1396_ ;
wire \myreg/_1397_ ;
wire \myreg/_1398_ ;
wire \myreg/_1399_ ;
wire \myreg/_1400_ ;
wire \myreg/_1401_ ;
wire \myreg/_1402_ ;
wire \myreg/_1403_ ;
wire \myreg/_1404_ ;
wire \myreg/_1405_ ;
wire \myreg/_1406_ ;
wire \myreg/_1407_ ;
wire \myreg/_1408_ ;
wire \myreg/_1409_ ;
wire \myreg/_1410_ ;
wire \myreg/_1411_ ;
wire \myreg/_1412_ ;
wire \myreg/_1413_ ;
wire \myreg/_1414_ ;
wire \myreg/_1415_ ;
wire \myreg/_1416_ ;
wire \myreg/_1417_ ;
wire \myreg/_1418_ ;
wire \myreg/_1419_ ;
wire \myreg/_1420_ ;
wire \myreg/_1421_ ;
wire \myreg/_1422_ ;
wire \myreg/_1423_ ;
wire \myreg/_1424_ ;
wire \myreg/_1425_ ;
wire \myreg/_1426_ ;
wire \myreg/_1427_ ;
wire \myreg/_1428_ ;
wire \myreg/_1429_ ;
wire \myreg/_1430_ ;
wire \myreg/_1431_ ;
wire \myreg/_1432_ ;
wire \myreg/_1433_ ;
wire \myreg/_1434_ ;
wire \myreg/_1435_ ;
wire \myreg/_1436_ ;
wire \myreg/_1437_ ;
wire \myreg/_1438_ ;
wire \myreg/_1439_ ;
wire \myreg/_1440_ ;
wire \myreg/_1441_ ;
wire \myreg/_1442_ ;
wire \myreg/_1443_ ;
wire \myreg/_1444_ ;
wire \myreg/_1445_ ;
wire \myreg/_1446_ ;
wire \myreg/_1447_ ;
wire \myreg/_1448_ ;
wire \myreg/_1449_ ;
wire \myreg/_1450_ ;
wire \myreg/_1451_ ;
wire \myreg/_1452_ ;
wire \myreg/_1453_ ;
wire \myreg/_1454_ ;
wire \myreg/_1455_ ;
wire \myreg/_1456_ ;
wire \myreg/_1457_ ;
wire \myreg/_1458_ ;
wire \myreg/_1459_ ;
wire \myreg/_1460_ ;
wire \myreg/_1461_ ;
wire \myreg/_1462_ ;
wire \myreg/_1463_ ;
wire \myreg/_1464_ ;
wire \myreg/_1465_ ;
wire \myreg/_1466_ ;
wire \myreg/_1467_ ;
wire \myreg/_1468_ ;
wire \myreg/_1469_ ;
wire \myreg/_1470_ ;
wire \myreg/_1471_ ;
wire \myreg/_1472_ ;
wire \myreg/_1473_ ;
wire \myreg/_1474_ ;
wire \myreg/_1475_ ;
wire \myreg/_1476_ ;
wire \myreg/_1477_ ;
wire \myreg/_1478_ ;
wire \myreg/_1479_ ;
wire \myreg/_1480_ ;
wire \myreg/_1481_ ;
wire \myreg/_1482_ ;
wire \myreg/_1483_ ;
wire \myreg/_1484_ ;
wire \myreg/_1485_ ;
wire \myreg/_1486_ ;
wire \myreg/_1487_ ;
wire \myreg/_1488_ ;
wire \myreg/_1489_ ;
wire \myreg/_1490_ ;
wire \myreg/_1491_ ;
wire \myreg/_1492_ ;
wire \myreg/_1493_ ;
wire \myreg/_1494_ ;
wire \myreg/_1495_ ;
wire \myreg/_1496_ ;
wire \myreg/_1497_ ;
wire \myreg/_1498_ ;
wire \myreg/_1499_ ;
wire \myreg/_1500_ ;
wire \myreg/_1501_ ;
wire \myreg/_1502_ ;
wire \myreg/_1503_ ;
wire \myreg/_1504_ ;
wire \myreg/_1505_ ;
wire \myreg/_1506_ ;
wire \myreg/_1507_ ;
wire \myreg/_1508_ ;
wire \myreg/_1509_ ;
wire \myreg/_1510_ ;
wire \myreg/_1511_ ;
wire \myreg/_1512_ ;
wire \myreg/_1513_ ;
wire \myreg/_1514_ ;
wire \myreg/_1515_ ;
wire \myreg/_1516_ ;
wire \myreg/_1517_ ;
wire \myreg/_1518_ ;
wire \myreg/_1519_ ;
wire \myreg/_1520_ ;
wire \myreg/_1521_ ;
wire \myreg/_1522_ ;
wire \myreg/_1523_ ;
wire \myreg/_1524_ ;
wire \myreg/_1525_ ;
wire \myreg/_1526_ ;
wire \myreg/_1527_ ;
wire \myreg/_1528_ ;
wire \myreg/_1529_ ;
wire \myreg/_1530_ ;
wire \myreg/_1531_ ;
wire \myreg/_1532_ ;
wire \myreg/_1533_ ;
wire \myreg/_1534_ ;
wire \myreg/_1535_ ;
wire \myreg/_1536_ ;
wire \myreg/_1537_ ;
wire \myreg/_1538_ ;
wire \myreg/_1539_ ;
wire \myreg/_1540_ ;
wire \myreg/_1541_ ;
wire \myreg/_1542_ ;
wire \myreg/_1543_ ;
wire \myreg/_1544_ ;
wire \myreg/_1545_ ;
wire \myreg/_1546_ ;
wire \myreg/_1547_ ;
wire \myreg/_1548_ ;
wire \myreg/_1549_ ;
wire \myreg/_1550_ ;
wire \myreg/_1551_ ;
wire \myreg/_1552_ ;
wire \myreg/_1553_ ;
wire \myreg/_1554_ ;
wire \myreg/_1555_ ;
wire \myreg/_1556_ ;
wire \myreg/_1557_ ;
wire \myreg/_1558_ ;
wire \myreg/_1559_ ;
wire \myreg/_1560_ ;
wire \myreg/_1561_ ;
wire \myreg/_1562_ ;
wire \myreg/_1563_ ;
wire \myreg/_1564_ ;
wire \myreg/_1565_ ;
wire \myreg/_1566_ ;
wire \myreg/_1567_ ;
wire \myreg/_1568_ ;
wire \myreg/_1569_ ;
wire \myreg/_1570_ ;
wire \myreg/_1571_ ;
wire \myreg/_1572_ ;
wire \myreg/_1573_ ;
wire \myreg/_1574_ ;
wire \myreg/_1575_ ;
wire \myreg/_1576_ ;
wire \myreg/_1577_ ;
wire \myreg/_1578_ ;
wire \myreg/_1579_ ;
wire \myreg/_1580_ ;
wire \myreg/_1581_ ;
wire \myreg/_1582_ ;
wire \myreg/_1583_ ;
wire \myreg/_1584_ ;
wire \myreg/_1585_ ;
wire \myreg/_1586_ ;
wire \myreg/_1587_ ;
wire \myreg/_1588_ ;
wire \myreg/_1589_ ;
wire \myreg/_1590_ ;
wire \myreg/_1591_ ;
wire \myreg/_1592_ ;
wire \myreg/_1593_ ;
wire \myreg/_1594_ ;
wire \myreg/_1595_ ;
wire \myreg/_1596_ ;
wire \myreg/_1597_ ;
wire \myreg/_1598_ ;
wire \myreg/_1599_ ;
wire \myreg/_1600_ ;
wire \myreg/_1601_ ;
wire \myreg/_1602_ ;
wire \myreg/_1603_ ;
wire \myreg/_1604_ ;
wire \myreg/_1605_ ;
wire \myreg/_1606_ ;
wire \myreg/_1607_ ;
wire \myreg/_1608_ ;
wire \myreg/_1609_ ;
wire \myreg/_1610_ ;
wire \myreg/_1611_ ;
wire \myreg/_1612_ ;
wire \myreg/_1613_ ;
wire \myreg/_1614_ ;
wire \myreg/_1615_ ;
wire \myreg/_1616_ ;
wire \myreg/_1617_ ;
wire \myreg/_1618_ ;
wire \myreg/_1619_ ;
wire \myreg/_1620_ ;
wire \myreg/_1621_ ;
wire \myreg/_1622_ ;
wire \myreg/_1623_ ;
wire \myreg/_1624_ ;
wire \myreg/_1625_ ;
wire \myreg/_1626_ ;
wire \myreg/_1627_ ;
wire \myreg/_1628_ ;
wire \myreg/_1629_ ;
wire \myreg/_1630_ ;
wire \myreg/_1631_ ;
wire \myreg/_1632_ ;
wire \myreg/_1633_ ;
wire \myreg/_1634_ ;
wire \myreg/_1635_ ;
wire \myreg/_1636_ ;
wire \myreg/_1637_ ;
wire \myreg/_1638_ ;
wire \myreg/_1639_ ;
wire \myreg/_1640_ ;
wire \myreg/_1641_ ;
wire \myreg/_1642_ ;
wire \myreg/_1643_ ;
wire \myreg/_1644_ ;
wire \myreg/_1645_ ;
wire \myreg/_1646_ ;
wire \myreg/_1647_ ;
wire \myreg/_1648_ ;
wire \myreg/_1649_ ;
wire \myreg/_1650_ ;
wire \myreg/_1651_ ;
wire \myreg/_1652_ ;
wire \myreg/_1653_ ;
wire \myreg/_1654_ ;
wire \myreg/_1655_ ;
wire \myreg/_1656_ ;
wire \myreg/_1657_ ;
wire \myreg/_1658_ ;
wire \myreg/_1659_ ;
wire \myreg/_1660_ ;
wire \myreg/_1661_ ;
wire \myreg/_1662_ ;
wire \myreg/_1663_ ;
wire \myreg/_1664_ ;
wire \myreg/_1665_ ;
wire \myreg/_1666_ ;
wire \myreg/_1667_ ;
wire \myreg/_1668_ ;
wire \myreg/_1669_ ;
wire \myreg/_1670_ ;
wire \myreg/_1671_ ;
wire \myreg/_1672_ ;
wire \myreg/_1673_ ;
wire \myreg/_1674_ ;
wire \myreg/_1675_ ;
wire \myreg/_1676_ ;
wire \myreg/_1677_ ;
wire \myreg/_1678_ ;
wire \myreg/_1679_ ;
wire \myreg/_1680_ ;
wire \myreg/_1681_ ;
wire \myreg/_1682_ ;
wire \myreg/_1683_ ;
wire \myreg/_1684_ ;
wire \myreg/_1685_ ;
wire \myreg/_1686_ ;
wire \myreg/_1687_ ;
wire \myreg/_1688_ ;
wire \myreg/_1689_ ;
wire \myreg/_1690_ ;
wire \myreg/_1691_ ;
wire \myreg/_1692_ ;
wire \myreg/_1693_ ;
wire \myreg/_1694_ ;
wire \myreg/_1695_ ;
wire \myreg/_1696_ ;
wire \myreg/_1697_ ;
wire \myreg/_1698_ ;
wire \myreg/_1699_ ;
wire \myreg/_1700_ ;
wire \myreg/_1701_ ;
wire \myreg/_1702_ ;
wire \myreg/_1703_ ;
wire \myreg/_1704_ ;
wire \myreg/_1705_ ;
wire \myreg/_1706_ ;
wire \myreg/_1707_ ;
wire \myreg/_1708_ ;
wire \myreg/_1709_ ;
wire \myreg/_1710_ ;
wire \myreg/_1711_ ;
wire \myreg/_1712_ ;
wire \myreg/_1713_ ;
wire \myreg/_1714_ ;
wire \myreg/_1715_ ;
wire \myreg/_1716_ ;
wire \myreg/_1717_ ;
wire \myreg/_1718_ ;
wire \myreg/_1719_ ;
wire \myreg/_1720_ ;
wire \myreg/_1721_ ;
wire \myreg/_1722_ ;
wire \myreg/_1723_ ;
wire \myreg/_1724_ ;
wire \myreg/_1725_ ;
wire \myreg/_1726_ ;
wire \myreg/_1727_ ;
wire \myreg/_1728_ ;
wire \myreg/_1729_ ;
wire \myreg/_1730_ ;
wire \myreg/_1731_ ;
wire \myreg/_1732_ ;
wire \myreg/_1733_ ;
wire \myreg/_1734_ ;
wire \myreg/_1735_ ;
wire \myreg/_1736_ ;
wire \myreg/_1737_ ;
wire \myreg/_1738_ ;
wire \myreg/_1739_ ;
wire \myreg/_1740_ ;
wire \myreg/_1741_ ;
wire \myreg/_1742_ ;
wire \myreg/_1743_ ;
wire \myreg/_1744_ ;
wire \myreg/_1745_ ;
wire \myreg/_1746_ ;
wire \myreg/_1747_ ;
wire \myreg/_1748_ ;
wire \myreg/_1749_ ;
wire \myreg/_1750_ ;
wire \myreg/_1751_ ;
wire \myreg/_1752_ ;
wire \myreg/_1753_ ;
wire \myreg/_1754_ ;
wire \myreg/_1755_ ;
wire \myreg/_1756_ ;
wire \myreg/_1757_ ;
wire \myreg/_1758_ ;
wire \myreg/_1759_ ;
wire \myreg/_1760_ ;
wire \myreg/_1761_ ;
wire \myreg/_1762_ ;
wire \myreg/_1763_ ;
wire \myreg/_1764_ ;
wire \myreg/_1765_ ;
wire \myreg/_1766_ ;
wire \myreg/_1767_ ;
wire \myreg/_1768_ ;
wire \myreg/_1769_ ;
wire \myreg/_1770_ ;
wire \myreg/_1771_ ;
wire \myreg/_1772_ ;
wire \myreg/_1773_ ;
wire \myreg/_1774_ ;
wire \myreg/_1775_ ;
wire \myreg/_1776_ ;
wire \myreg/_1777_ ;
wire \myreg/_1778_ ;
wire \myreg/_1779_ ;
wire \myreg/_1780_ ;
wire \myreg/_1781_ ;
wire \myreg/_1782_ ;
wire \myreg/_1783_ ;
wire \myreg/_1784_ ;
wire \myreg/_1785_ ;
wire \myreg/_1786_ ;
wire \myreg/_1787_ ;
wire \myreg/_1788_ ;
wire \myreg/_1789_ ;
wire \myreg/_1790_ ;
wire \myreg/_1791_ ;
wire \myreg/_1792_ ;
wire \myreg/_1793_ ;
wire \myreg/_1794_ ;
wire \myreg/_1795_ ;
wire \myreg/_1796_ ;
wire \myreg/_1797_ ;
wire \myreg/_1798_ ;
wire \myreg/_1799_ ;
wire \myreg/_1800_ ;
wire \myreg/_1801_ ;
wire \myreg/_1802_ ;
wire \myreg/_1803_ ;
wire \myreg/_1804_ ;
wire \myreg/_1805_ ;
wire \myreg/_1806_ ;
wire \myreg/_1807_ ;
wire \myreg/_1808_ ;
wire \myreg/_1809_ ;
wire \myreg/_1810_ ;
wire \myreg/_1811_ ;
wire \myreg/_1812_ ;
wire \myreg/_1813_ ;
wire \myreg/_1814_ ;
wire \myreg/_1815_ ;
wire \myreg/_1816_ ;
wire \myreg/_1817_ ;
wire \myreg/_1818_ ;
wire \myreg/_1819_ ;
wire \myreg/_1820_ ;
wire \myreg/_1821_ ;
wire \myreg/_1822_ ;
wire \myreg/_1823_ ;
wire \myreg/_1824_ ;
wire \myreg/_1825_ ;
wire \myreg/_1826_ ;
wire \myreg/_1827_ ;
wire \myreg/_1828_ ;
wire \myreg/_1829_ ;
wire \myreg/_1830_ ;
wire \myreg/_1831_ ;
wire \myreg/_1832_ ;
wire \myreg/_1833_ ;
wire \myreg/_1834_ ;
wire \myreg/_1835_ ;
wire \myreg/_1836_ ;
wire \myreg/_1837_ ;
wire \myreg/_1838_ ;
wire \myreg/_1839_ ;
wire \myreg/_1840_ ;
wire \myreg/_1841_ ;
wire \myreg/_1842_ ;
wire \myreg/_1843_ ;
wire \myreg/_1844_ ;
wire \myreg/_1845_ ;
wire \myreg/_1846_ ;
wire \myreg/_1847_ ;
wire \myreg/_1848_ ;
wire \myreg/_1849_ ;
wire \myreg/_1850_ ;
wire \myreg/_1851_ ;
wire \myreg/_1852_ ;
wire \myreg/_1853_ ;
wire \myreg/_1854_ ;
wire \myreg/_1855_ ;
wire \myreg/_1856_ ;
wire \myreg/_1857_ ;
wire \myreg/_1858_ ;
wire \myreg/_1859_ ;
wire \myreg/_1860_ ;
wire \myreg/_1861_ ;
wire \myreg/_1862_ ;
wire \myreg/_1863_ ;
wire \myreg/_1864_ ;
wire \myreg/_1865_ ;
wire \myreg/_1866_ ;
wire \myreg/_1867_ ;
wire \myreg/_1868_ ;
wire \myreg/_1869_ ;
wire \myreg/_1870_ ;
wire \myreg/_1871_ ;
wire \myreg/_1872_ ;
wire \myreg/_1873_ ;
wire \myreg/_1874_ ;
wire \myreg/_1875_ ;
wire \myreg/_1876_ ;
wire \myreg/_1877_ ;
wire \myreg/_1878_ ;
wire \myreg/_1879_ ;
wire \myreg/_1880_ ;
wire \myreg/_1881_ ;
wire \myreg/_1882_ ;
wire \myreg/_1883_ ;
wire \myreg/_1884_ ;
wire \myreg/_1885_ ;
wire \myreg/_1886_ ;
wire \myreg/_1887_ ;
wire \myreg/_1888_ ;
wire \myreg/_1889_ ;
wire \myreg/_1890_ ;
wire \myreg/_1891_ ;
wire \myreg/_1892_ ;
wire \myreg/_1893_ ;
wire \myreg/_1894_ ;
wire \myreg/_1895_ ;
wire \myreg/_1896_ ;
wire \myreg/_1897_ ;
wire \myreg/_1898_ ;
wire \myreg/_1899_ ;
wire \myreg/_1900_ ;
wire \myreg/_1901_ ;
wire \myreg/_1902_ ;
wire \myreg/_1903_ ;
wire \myreg/_1904_ ;
wire \myreg/_1905_ ;
wire \myreg/_1906_ ;
wire \myreg/_1907_ ;
wire \myreg/_1908_ ;
wire \myreg/_1909_ ;
wire \myreg/_1910_ ;
wire \myreg/_1911_ ;
wire \myreg/_1912_ ;
wire \myreg/_1913_ ;
wire \myreg/_1914_ ;
wire \myreg/_1915_ ;
wire \myreg/_1916_ ;
wire \myreg/_1917_ ;
wire \myreg/_1918_ ;
wire \myreg/_1919_ ;
wire \myreg/_1920_ ;
wire \myreg/_1921_ ;
wire \myreg/_1922_ ;
wire \myreg/_1923_ ;
wire \myreg/_1924_ ;
wire \myreg/_1925_ ;
wire \myreg/_1926_ ;
wire \myreg/_1927_ ;
wire \myreg/_1928_ ;
wire \myreg/_1929_ ;
wire \myreg/_1930_ ;
wire \myreg/_1931_ ;
wire \myreg/_1932_ ;
wire \myreg/_1933_ ;
wire \myreg/_1934_ ;
wire \myreg/_1935_ ;
wire \myreg/_1936_ ;
wire \myreg/_1937_ ;
wire \myreg/_1938_ ;
wire \myreg/_1939_ ;
wire \myreg/_1940_ ;
wire \myreg/_1941_ ;
wire \myreg/_1942_ ;
wire \myreg/_1943_ ;
wire \myreg/_1944_ ;
wire \myreg/_1945_ ;
wire \myreg/_1946_ ;
wire \myreg/_1947_ ;
wire \myreg/_1948_ ;
wire \myreg/_1949_ ;
wire \myreg/_1950_ ;
wire \myreg/_1951_ ;
wire \myreg/_1952_ ;
wire \myreg/_1953_ ;
wire \myreg/_1954_ ;
wire \myreg/_1955_ ;
wire \myreg/_1956_ ;
wire \myreg/_1957_ ;
wire \myreg/_1958_ ;
wire \myreg/_1959_ ;
wire \myreg/_1960_ ;
wire \myreg/_1961_ ;
wire \myreg/_1962_ ;
wire \myreg/_1963_ ;
wire \myreg/_1964_ ;
wire \myreg/_1965_ ;
wire \myreg/_1966_ ;
wire \myreg/_1967_ ;
wire \myreg/_1968_ ;
wire \myreg/_1969_ ;
wire \myreg/_1970_ ;
wire \myreg/_1971_ ;
wire \myreg/_1972_ ;
wire \myreg/_1973_ ;
wire \myreg/_1974_ ;
wire \myreg/_1975_ ;
wire \myreg/_1976_ ;
wire \myreg/_1977_ ;
wire \myreg/_1978_ ;
wire \myreg/_1979_ ;
wire \myreg/_1980_ ;
wire \myreg/_1981_ ;
wire \myreg/_1982_ ;
wire \myreg/_1983_ ;
wire \myreg/_1984_ ;
wire \myreg/_1985_ ;
wire \myreg/_1986_ ;
wire \myreg/_1987_ ;
wire \myreg/_1988_ ;
wire \myreg/_1989_ ;
wire \myreg/_1990_ ;
wire \myreg/_1991_ ;
wire \myreg/_1992_ ;
wire \myreg/_1993_ ;
wire \myreg/_1994_ ;
wire \myreg/_1995_ ;
wire \myreg/_1996_ ;
wire \myreg/_1997_ ;
wire \myreg/_1998_ ;
wire \myreg/_1999_ ;
wire \myreg/_2000_ ;
wire \myreg/_2001_ ;
wire \myreg/_2002_ ;
wire \myreg/_2003_ ;
wire \myreg/_2004_ ;
wire \myreg/_2005_ ;
wire \myreg/_2006_ ;
wire \myreg/_2007_ ;
wire \myreg/_2008_ ;
wire \myreg/_2009_ ;
wire \myreg/_2010_ ;
wire \myreg/_2011_ ;
wire \myreg/_2012_ ;
wire \myreg/_2013_ ;
wire \myreg/_2014_ ;
wire \myreg/_2015_ ;
wire \myreg/_2016_ ;
wire \myreg/_2017_ ;
wire \myreg/_2018_ ;
wire \myreg/_2019_ ;
wire \myreg/_2020_ ;
wire \myreg/_2021_ ;
wire \myreg/_2022_ ;
wire \myreg/_2023_ ;
wire \myreg/_2024_ ;
wire \myreg/_2025_ ;
wire \myreg/_2026_ ;
wire \myreg/_2027_ ;
wire \myreg/_2028_ ;
wire \myreg/_2029_ ;
wire \myreg/_2030_ ;
wire \myreg/_2031_ ;
wire \myreg/_2032_ ;
wire \myreg/_2033_ ;
wire \myreg/_2034_ ;
wire \myreg/_2035_ ;
wire \myreg/_2036_ ;
wire \myreg/_2037_ ;
wire \myreg/_2038_ ;
wire \myreg/_2039_ ;
wire \myreg/_2040_ ;
wire \myreg/_2041_ ;
wire \myreg/_2042_ ;
wire \myreg/_2043_ ;
wire \myreg/_2044_ ;
wire \myreg/_2045_ ;
wire \myreg/_2046_ ;
wire \myreg/_2047_ ;
wire \myreg/_2048_ ;
wire \myreg/_2049_ ;
wire \myreg/_2050_ ;
wire \myreg/_2051_ ;
wire \myreg/_2052_ ;
wire \myreg/_2053_ ;
wire \myreg/_2054_ ;
wire \myreg/_2055_ ;
wire \myreg/_2056_ ;
wire \myreg/_2057_ ;
wire \myreg/_2058_ ;
wire \myreg/_2059_ ;
wire \myreg/_2060_ ;
wire \myreg/_2061_ ;
wire \myreg/_2062_ ;
wire \myreg/_2063_ ;
wire \myreg/_2064_ ;
wire \myreg/_2065_ ;
wire \myreg/_2066_ ;
wire \myreg/_2067_ ;
wire \myreg/_2068_ ;
wire \myreg/_2069_ ;
wire \myreg/_2070_ ;
wire \myreg/_2071_ ;
wire \myreg/_2072_ ;
wire \myreg/_2073_ ;
wire \myreg/_2074_ ;
wire \myreg/_2075_ ;
wire \myreg/_2076_ ;
wire \myreg/_2077_ ;
wire \myreg/_2078_ ;
wire \myreg/_2079_ ;
wire \myreg/_2080_ ;
wire \myreg/_2081_ ;
wire \myreg/_2082_ ;
wire \myreg/_2083_ ;
wire \myreg/_2084_ ;
wire \myreg/_2085_ ;
wire \myreg/_2086_ ;
wire \myreg/_2087_ ;
wire \myreg/_2088_ ;
wire \myreg/_2089_ ;
wire \myreg/_2090_ ;
wire \myreg/_2091_ ;
wire \myreg/_2092_ ;
wire \myreg/_2093_ ;
wire \myreg/_2094_ ;
wire \myreg/_2095_ ;
wire \myreg/_2096_ ;
wire \myreg/_2097_ ;
wire \myreg/_2098_ ;
wire \myreg/_2099_ ;
wire \myreg/_2100_ ;
wire \myreg/_2101_ ;
wire \myreg/_2102_ ;
wire \myreg/_2103_ ;
wire \myreg/_2104_ ;
wire \myreg/_2105_ ;
wire \myreg/_2106_ ;
wire \myreg/_2107_ ;
wire \myreg/_2108_ ;
wire \myreg/_2109_ ;
wire \myreg/_2110_ ;
wire \myreg/_2111_ ;
wire \myreg/_2112_ ;
wire \myreg/_2113_ ;
wire \myreg/_2114_ ;
wire \myreg/_2115_ ;
wire \myreg/_2116_ ;
wire \myreg/_2117_ ;
wire \myreg/_2118_ ;
wire \myreg/_2119_ ;
wire \myreg/_2120_ ;
wire \myreg/_2121_ ;
wire \myreg/_2122_ ;
wire \myreg/_2123_ ;
wire \myreg/_2124_ ;
wire \myreg/_2125_ ;
wire \myreg/_2126_ ;
wire \myreg/_2127_ ;
wire \myreg/_2128_ ;
wire \myreg/_2129_ ;
wire \myreg/_2130_ ;
wire \myreg/_2131_ ;
wire \myreg/_2132_ ;
wire \myreg/_2133_ ;
wire \myreg/_2134_ ;
wire \myreg/_2135_ ;
wire \myreg/_2136_ ;
wire \myreg/_2137_ ;
wire \myreg/_2138_ ;
wire \myreg/_2139_ ;
wire \myreg/_2140_ ;
wire \myreg/_2141_ ;
wire \myreg/_2142_ ;
wire \myreg/_2143_ ;
wire \myreg/_2144_ ;
wire \myreg/_2145_ ;
wire \myreg/_2146_ ;
wire \myreg/_2147_ ;
wire \myreg/_2148_ ;
wire \myreg/_2149_ ;
wire \myreg/_2150_ ;
wire \myreg/_2151_ ;
wire \myreg/_2152_ ;
wire \myreg/_2153_ ;
wire \myreg/_2154_ ;
wire \myreg/_2155_ ;
wire \myreg/_2156_ ;
wire \myreg/_2157_ ;
wire \myreg/_2158_ ;
wire \myreg/_2159_ ;
wire \myreg/_2160_ ;
wire \myreg/_2161_ ;
wire \myreg/_2162_ ;
wire \myreg/_2163_ ;
wire \myreg/_2164_ ;
wire \myreg/_2165_ ;
wire \myreg/_2166_ ;
wire \myreg/_2167_ ;
wire \myreg/_2168_ ;
wire \myreg/_2169_ ;
wire \myreg/_2170_ ;
wire \myreg/_2171_ ;
wire \myreg/_2172_ ;
wire \myreg/_2173_ ;
wire \myreg/_2174_ ;
wire \myreg/_2175_ ;
wire \myreg/_2176_ ;
wire \myreg/_2177_ ;
wire \myreg/_2178_ ;
wire \myreg/_2179_ ;
wire \myreg/_2180_ ;
wire \myreg/_2181_ ;
wire \myreg/_2182_ ;
wire \myreg/_2183_ ;
wire \myreg/_2184_ ;
wire \myreg/_2185_ ;
wire \myreg/_2186_ ;
wire \myreg/_2187_ ;
wire \myreg/_2188_ ;
wire \myreg/_2189_ ;
wire \myreg/_2190_ ;
wire \myreg/_2191_ ;
wire \myreg/_2192_ ;
wire \myreg/_2193_ ;
wire \myreg/_2194_ ;
wire \myreg/_2195_ ;
wire \myreg/_2196_ ;
wire \myreg/_2197_ ;
wire \myreg/_2198_ ;
wire \myreg/_2199_ ;
wire \myreg/_2200_ ;
wire \myreg/_2201_ ;
wire \myreg/_2202_ ;
wire \myreg/_2203_ ;
wire \myreg/_2204_ ;
wire \myreg/_2205_ ;
wire \myreg/_2206_ ;
wire \myreg/_2207_ ;
wire \myreg/_2208_ ;
wire \myreg/_2209_ ;
wire \myreg/_2210_ ;
wire \myreg/_2211_ ;
wire \myreg/_2212_ ;
wire \myreg/_2213_ ;
wire \myreg/_2214_ ;
wire \myreg/_2215_ ;
wire \myreg/_2216_ ;
wire \myreg/_2217_ ;
wire \myreg/_2218_ ;
wire \myreg/_2219_ ;
wire \myreg/_2220_ ;
wire \myreg/_2221_ ;
wire \myreg/_2222_ ;
wire \myreg/_2223_ ;
wire \myreg/_2224_ ;
wire \myreg/_2225_ ;
wire \myreg/_2226_ ;
wire \myreg/_2227_ ;
wire \myreg/_2228_ ;
wire \myreg/_2229_ ;
wire \myreg/_2230_ ;
wire \myreg/_2231_ ;
wire \myreg/_2232_ ;
wire \myreg/_2233_ ;
wire \myreg/_2234_ ;
wire \myreg/_2235_ ;
wire \myreg/_2236_ ;
wire \myreg/_2237_ ;
wire \myreg/_2238_ ;
wire \myreg/_2239_ ;
wire \myreg/_2240_ ;
wire \myreg/_2241_ ;
wire \myreg/_2242_ ;
wire \myreg/_2243_ ;
wire \myreg/_2244_ ;
wire \myreg/_2245_ ;
wire \myreg/_2246_ ;
wire \myreg/_2247_ ;
wire \myreg/_2248_ ;
wire \myreg/_2249_ ;
wire \myreg/_2250_ ;
wire \myreg/_2251_ ;
wire \myreg/_2252_ ;
wire \myreg/_2253_ ;
wire \myreg/_2254_ ;
wire \myreg/_2255_ ;
wire \myreg/_2256_ ;
wire \myreg/_2257_ ;
wire \myreg/_2258_ ;
wire \myreg/_2259_ ;
wire \myreg/_2260_ ;
wire \myreg/_2261_ ;
wire \myreg/_2262_ ;
wire \myreg/_2263_ ;
wire \myreg/_2264_ ;
wire \myreg/_2265_ ;
wire \myreg/_2266_ ;
wire \myreg/_2267_ ;
wire \myreg/_2268_ ;
wire \myreg/_2269_ ;
wire \myreg/_2270_ ;
wire \myreg/_2271_ ;
wire \myreg/_2272_ ;
wire \myreg/_2273_ ;
wire \myreg/_2274_ ;
wire \myreg/_2275_ ;
wire \myreg/_2276_ ;
wire \myreg/_2277_ ;
wire \myreg/_2278_ ;
wire \myreg/_2279_ ;
wire \myreg/_2280_ ;
wire \myreg/_2281_ ;
wire \myreg/_2282_ ;
wire \myreg/_2283_ ;
wire \myreg/_2284_ ;
wire \myreg/_2285_ ;
wire \myreg/_2286_ ;
wire \myreg/_2287_ ;
wire \myreg/_2288_ ;
wire \myreg/_2289_ ;
wire \myreg/_2290_ ;
wire \myreg/_2291_ ;
wire \myreg/_2292_ ;
wire \myreg/_2293_ ;
wire \myreg/_2294_ ;
wire \myreg/_2295_ ;
wire \myreg/_2296_ ;
wire \myreg/_2297_ ;
wire \myreg/_2298_ ;
wire \myreg/_2299_ ;
wire \myreg/_2300_ ;
wire \myreg/_2301_ ;
wire \myreg/_2302_ ;
wire \myreg/_2303_ ;
wire \myreg/_2304_ ;
wire \myreg/_2305_ ;
wire \myreg/_2306_ ;
wire \myreg/_2307_ ;
wire \myreg/_2308_ ;
wire \myreg/_2309_ ;
wire \myreg/_2310_ ;
wire \myreg/_2311_ ;
wire \myreg/_2312_ ;
wire \myreg/_2313_ ;
wire \myreg/_2314_ ;
wire \myreg/_2315_ ;
wire \myreg/_2316_ ;
wire \myreg/_2317_ ;
wire \myreg/_2318_ ;
wire \myreg/_2319_ ;
wire \myreg/_2320_ ;
wire \myreg/_2321_ ;
wire \myreg/_2322_ ;
wire \myreg/_2323_ ;
wire \myreg/_2324_ ;
wire \myreg/_2325_ ;
wire \myreg/_2326_ ;
wire \myreg/_2327_ ;
wire \myreg/_2328_ ;
wire \myreg/_2329_ ;
wire \myreg/_2330_ ;
wire \myreg/_2331_ ;
wire \myreg/_2332_ ;
wire \myreg/_2333_ ;
wire \myreg/_2334_ ;
wire \myreg/_2335_ ;
wire \myreg/_2336_ ;
wire \myreg/_2337_ ;
wire \myreg/_2338_ ;
wire \myreg/_2339_ ;
wire \myreg/_2340_ ;
wire \myreg/_2341_ ;
wire \myreg/_2342_ ;
wire \myreg/_2343_ ;
wire \myreg/_2344_ ;
wire \myreg/_2345_ ;
wire \myreg/_2346_ ;
wire \myreg/_2347_ ;
wire \myreg/_2348_ ;
wire \myreg/_2349_ ;
wire \myreg/_2350_ ;
wire \myreg/_2351_ ;
wire \myreg/_2352_ ;
wire \myreg/_2353_ ;
wire \myreg/_2354_ ;
wire \myreg/_2355_ ;
wire \myreg/_2356_ ;
wire \myreg/_2357_ ;
wire \myreg/_2358_ ;
wire \myreg/_2359_ ;
wire \myreg/_2360_ ;
wire \myreg/_2361_ ;
wire \myreg/_2362_ ;
wire \myreg/_2363_ ;
wire \myreg/_2364_ ;
wire \myreg/_2365_ ;
wire \myreg/_2366_ ;
wire \myreg/_2367_ ;
wire \myreg/_2368_ ;
wire \myreg/_2369_ ;
wire \myreg/_2370_ ;
wire \myreg/_2371_ ;
wire \myreg/_2372_ ;
wire \myreg/_2373_ ;
wire \myreg/_2374_ ;
wire \myreg/_2375_ ;
wire \myreg/_2376_ ;
wire \myreg/_2377_ ;
wire \myreg/_2378_ ;
wire \myreg/_2379_ ;
wire \myreg/_2380_ ;
wire \myreg/_2381_ ;
wire \myreg/_2382_ ;
wire \myreg/_2383_ ;
wire \myreg/_2384_ ;
wire \myreg/_2385_ ;
wire \myreg/_2386_ ;
wire \myreg/_2387_ ;
wire \myreg/_2388_ ;
wire \myreg/_2389_ ;
wire \myreg/_2390_ ;
wire \myreg/_2391_ ;
wire \myreg/_2392_ ;
wire \myreg/_2393_ ;
wire \myreg/_2394_ ;
wire \myreg/_2395_ ;
wire \myreg/_2396_ ;
wire \myreg/_2397_ ;
wire \myreg/_2398_ ;
wire \myreg/_2399_ ;
wire \myreg/_2400_ ;
wire \myreg/_2401_ ;
wire \myreg/_2402_ ;
wire \myreg/_2403_ ;
wire \myreg/_2404_ ;
wire \myreg/_2405_ ;
wire \myreg/_2406_ ;
wire \myreg/_2407_ ;
wire \myreg/_2408_ ;
wire \myreg/_2409_ ;
wire \myreg/_2410_ ;
wire \myreg/_2411_ ;
wire \myreg/_2412_ ;
wire \myreg/_2413_ ;
wire \myreg/_2414_ ;
wire \myreg/_2415_ ;
wire \myreg/_2416_ ;
wire \myreg/_2417_ ;
wire \myreg/_2418_ ;
wire \myreg/_2419_ ;
wire \myreg/_2420_ ;
wire \myreg/_2421_ ;
wire \myreg/_2422_ ;
wire \myreg/_2423_ ;
wire \myreg/_2424_ ;
wire \myreg/_2425_ ;
wire \myreg/_2426_ ;
wire \myreg/_2427_ ;
wire \myreg/_2428_ ;
wire \myreg/_2429_ ;
wire \myreg/_2430_ ;
wire \myreg/_2431_ ;
wire \myreg/_2432_ ;
wire \myreg/_2433_ ;
wire \myreg/_2434_ ;
wire \myreg/_2435_ ;
wire \myreg/_2436_ ;
wire \myreg/_2437_ ;
wire \myreg/_2438_ ;
wire \myreg/_2439_ ;
wire \myreg/_2440_ ;
wire \myreg/_2441_ ;
wire \myreg/_2442_ ;
wire \myreg/_2443_ ;
wire \myreg/_2444_ ;
wire \myreg/_2445_ ;
wire \myreg/_2446_ ;
wire \myreg/_2447_ ;
wire \myreg/_2448_ ;
wire \myreg/_2449_ ;
wire \myreg/_2450_ ;
wire \myreg/_2451_ ;
wire \myreg/_2452_ ;
wire \myreg/_2453_ ;
wire \myreg/_2454_ ;
wire \myreg/_2455_ ;
wire \myreg/_2456_ ;
wire \myreg/_2457_ ;
wire \myreg/_2458_ ;
wire \myreg/_2459_ ;
wire \myreg/_2460_ ;
wire \myreg/_2461_ ;
wire \myreg/_2462_ ;
wire \myreg/_2463_ ;
wire \myreg/_2464_ ;
wire \myreg/_2465_ ;
wire \myreg/_2466_ ;
wire \myreg/_2467_ ;
wire \myreg/_2468_ ;
wire \myreg/_2469_ ;
wire \myreg/_2470_ ;
wire \myreg/_2471_ ;
wire \myreg/_2472_ ;
wire \myreg/_2473_ ;
wire \myreg/_2474_ ;
wire \myreg/_2475_ ;
wire \myreg/_2476_ ;
wire \myreg/_2477_ ;
wire \myreg/_2478_ ;
wire \myreg/_2479_ ;
wire \myreg/_2480_ ;
wire \myreg/_2481_ ;
wire \myreg/_2482_ ;
wire \myreg/_2483_ ;
wire \myreg/_2484_ ;
wire \myreg/_2485_ ;
wire \myreg/_2486_ ;
wire \myreg/_2487_ ;
wire \myreg/_2488_ ;
wire \myreg/_2489_ ;
wire \myreg/_2490_ ;
wire \myreg/_2491_ ;
wire \myreg/_2492_ ;
wire \myreg/_2493_ ;
wire \myreg/_2494_ ;
wire \myreg/_2495_ ;
wire \myreg/_2496_ ;
wire \myreg/_2497_ ;
wire \myreg/_2498_ ;
wire \myreg/_2499_ ;
wire \myreg/_2500_ ;
wire \myreg/_2501_ ;
wire \myreg/_2502_ ;
wire \myreg/_2503_ ;
wire \myreg/_2504_ ;
wire \myreg/_2505_ ;
wire \myreg/_2506_ ;
wire \myreg/_2507_ ;
wire \myreg/_2508_ ;
wire \myreg/_2509_ ;
wire \myreg/_2510_ ;
wire \myreg/_2511_ ;
wire \myreg/_2512_ ;
wire \myreg/_2513_ ;
wire \myreg/_2514_ ;
wire \myreg/_2515_ ;
wire \myreg/_2516_ ;
wire \myreg/_2517_ ;
wire \myreg/_2518_ ;
wire \myreg/_2519_ ;
wire \myreg/_2520_ ;
wire \myreg/_2521_ ;
wire \myreg/_2522_ ;
wire \myreg/_2523_ ;
wire \myreg/_2524_ ;
wire \myreg/_2525_ ;
wire \myreg/_2526_ ;
wire \myreg/_2527_ ;
wire \myreg/_2528_ ;
wire \myreg/_2529_ ;
wire \myreg/_2530_ ;
wire \myreg/_2531_ ;
wire \myreg/_2532_ ;
wire \myreg/_2533_ ;
wire \myreg/_2534_ ;
wire \myreg/_2535_ ;
wire \myreg/_2536_ ;
wire \myreg/_2537_ ;
wire \myreg/_2538_ ;
wire \myreg/_2539_ ;
wire \myreg/_2540_ ;
wire \myreg/_2541_ ;
wire \myreg/_2542_ ;
wire \myreg/_2543_ ;
wire \myreg/_2544_ ;
wire \myreg/_2545_ ;
wire \myreg/_2546_ ;
wire \myreg/_2547_ ;
wire \myreg/_2548_ ;
wire \myreg/_2549_ ;
wire \myreg/_2550_ ;
wire \myreg/_2551_ ;
wire \myreg/_2552_ ;
wire \myreg/_2553_ ;
wire \myreg/_2554_ ;
wire \myreg/_2555_ ;
wire \myreg/_2556_ ;
wire \myreg/_2557_ ;
wire \myreg/_2558_ ;
wire \myreg/_2559_ ;
wire \myreg/_2560_ ;
wire \myreg/_2561_ ;
wire \myreg/_2562_ ;
wire \myreg/_2563_ ;
wire \myreg/_2564_ ;
wire \myreg/_2565_ ;
wire \myreg/_2566_ ;
wire \myreg/_2567_ ;
wire \myreg/_2568_ ;
wire \myreg/_2569_ ;
wire \myreg/_2570_ ;
wire \myreg/_2571_ ;
wire \myreg/_2572_ ;
wire \myreg/_2573_ ;
wire \myreg/_2574_ ;
wire \myreg/_2575_ ;
wire \myreg/_2576_ ;
wire \myreg/_2577_ ;
wire \myreg/_2578_ ;
wire \myreg/_2579_ ;
wire \myreg/_2580_ ;
wire \myreg/_2581_ ;
wire \myreg/_2582_ ;
wire \myreg/_2583_ ;
wire \myreg/_2584_ ;
wire \myreg/_2585_ ;
wire \myreg/_2586_ ;
wire \myreg/_2587_ ;
wire \myreg/_2588_ ;
wire \myreg/_2589_ ;
wire \myreg/_2590_ ;
wire \myreg/_2591_ ;
wire \myreg/_2592_ ;
wire \myreg/_2593_ ;
wire \myreg/_2594_ ;
wire \myreg/_2595_ ;
wire \myreg/_2596_ ;
wire \myreg/_2597_ ;
wire \myreg/_2598_ ;
wire \myreg/_2599_ ;
wire \myreg/_2600_ ;
wire \myreg/_2601_ ;
wire \myreg/_2602_ ;
wire \myreg/_2603_ ;
wire \myreg/_2604_ ;
wire \myreg/_2605_ ;
wire \myreg/_2606_ ;
wire \myreg/_2607_ ;
wire \myreg/_2608_ ;
wire \myreg/_2609_ ;
wire \myreg/_2610_ ;
wire \myreg/_2611_ ;
wire \myreg/_2612_ ;
wire \myreg/_2613_ ;
wire \myreg/_2614_ ;
wire \myreg/_2615_ ;
wire \myreg/_2616_ ;
wire \myreg/_2617_ ;
wire \myreg/_2618_ ;
wire \myreg/_2619_ ;
wire \myreg/_2620_ ;
wire \myreg/_2621_ ;
wire \myreg/_2622_ ;
wire \myreg/_2623_ ;
wire \myreg/_2624_ ;
wire \myreg/_2625_ ;
wire \myreg/_2626_ ;
wire \myreg/_2627_ ;
wire \myreg/_2628_ ;
wire \myreg/_2629_ ;
wire \myreg/_2630_ ;
wire \myreg/_2631_ ;
wire \myreg/_2632_ ;
wire \myreg/_2633_ ;
wire \myreg/_2634_ ;
wire \myreg/_2635_ ;
wire \myreg/_2636_ ;
wire \myreg/_2637_ ;
wire \myreg/_2638_ ;
wire \myreg/_2639_ ;
wire \myreg/_2640_ ;
wire \myreg/_2641_ ;
wire \myreg/_2642_ ;
wire \myreg/_2643_ ;
wire \myreg/_2644_ ;
wire \myreg/_2645_ ;
wire \myreg/_2646_ ;
wire \myreg/_2647_ ;
wire \myreg/_2648_ ;
wire \myreg/_2649_ ;
wire \myreg/_2650_ ;
wire \myreg/_2651_ ;
wire \myreg/_2652_ ;
wire \myreg/_2653_ ;
wire \myreg/_2654_ ;
wire \myreg/_2655_ ;
wire \myreg/_2656_ ;
wire \myreg/_2657_ ;
wire \myreg/_2658_ ;
wire \myreg/_2659_ ;
wire \myreg/_2660_ ;
wire \myreg/_2661_ ;
wire \myreg/_2662_ ;
wire \myreg/_2663_ ;
wire \myreg/_2664_ ;
wire \myreg/_2665_ ;
wire \myreg/_2666_ ;
wire \myreg/_2667_ ;
wire \myreg/_2668_ ;
wire \myreg/_2669_ ;
wire \myreg/_2670_ ;
wire \myreg/_2671_ ;
wire \myreg/_2672_ ;
wire \myreg/_2673_ ;
wire \myreg/_2674_ ;
wire \myreg/_2675_ ;
wire \myreg/_2676_ ;
wire \myreg/_2677_ ;
wire \myreg/_2678_ ;
wire \myreg/_2679_ ;
wire \myreg/_2680_ ;
wire \myreg/_2681_ ;
wire \myreg/_2682_ ;
wire \myreg/_2683_ ;
wire \myreg/_2684_ ;
wire \myreg/_2685_ ;
wire \myreg/_2686_ ;
wire \myreg/_2687_ ;
wire \myreg/_2688_ ;
wire \myreg/_2689_ ;
wire \myreg/_2690_ ;
wire \myreg/_2691_ ;
wire \myreg/_2692_ ;
wire \myreg/_2693_ ;
wire \myreg/_2694_ ;
wire \myreg/_2695_ ;
wire \myreg/_2696_ ;
wire \myreg/_2697_ ;
wire \myreg/_2698_ ;
wire \myreg/_2699_ ;
wire \myreg/_2700_ ;
wire \myreg/_2701_ ;
wire \myreg/_2702_ ;
wire \myreg/_2703_ ;
wire \myreg/_2704_ ;
wire \myreg/_2705_ ;
wire \myreg/_2706_ ;
wire \myreg/_2707_ ;
wire \myreg/_2708_ ;
wire \myreg/_2709_ ;
wire \myreg/_2710_ ;
wire \myreg/_2711_ ;
wire \myreg/_2712_ ;
wire \myreg/_2713_ ;
wire \myreg/_2714_ ;
wire \myreg/_2715_ ;
wire \myreg/_2716_ ;
wire \myreg/_2717_ ;
wire \myreg/_2718_ ;
wire \myreg/_2719_ ;
wire \myreg/_2720_ ;
wire \myreg/_2721_ ;
wire \myreg/_2722_ ;
wire \myreg/_2723_ ;
wire \myreg/_2724_ ;
wire \myreg/_2725_ ;
wire \myreg/_2726_ ;
wire \myreg/_2727_ ;
wire \myreg/_2728_ ;
wire \myreg/_2729_ ;
wire \myreg/_2730_ ;
wire \myreg/_2731_ ;
wire \myreg/_2732_ ;
wire \myreg/_2733_ ;
wire \myreg/_2734_ ;
wire \myreg/_2735_ ;
wire \myreg/_2736_ ;
wire \myreg/_2737_ ;
wire \myreg/_2738_ ;
wire \myreg/_2739_ ;
wire \myreg/_2740_ ;
wire \myreg/_2741_ ;
wire \myreg/_2742_ ;
wire \myreg/_2743_ ;
wire \myreg/_2744_ ;
wire \myreg/_2745_ ;
wire \myreg/_2746_ ;
wire \myreg/_2747_ ;
wire \myreg/_2748_ ;
wire \myreg/_2749_ ;
wire \myreg/_2750_ ;
wire \myreg/_2751_ ;
wire \myreg/_2752_ ;
wire \myreg/_2753_ ;
wire \myreg/_2754_ ;
wire \myreg/_2755_ ;
wire \myreg/_2756_ ;
wire \myreg/_2757_ ;
wire \myreg/_2758_ ;
wire \myreg/_2759_ ;
wire \myreg/_2760_ ;
wire \myreg/_2761_ ;
wire \myreg/_2762_ ;
wire \myreg/_2763_ ;
wire \myreg/_2764_ ;
wire \myreg/_2765_ ;
wire \myreg/_2766_ ;
wire \myreg/_2767_ ;
wire \myreg/_2768_ ;
wire \myreg/_2769_ ;
wire \myreg/_2770_ ;
wire \myreg/_2771_ ;
wire \myreg/_2772_ ;
wire \myreg/_2773_ ;
wire \myreg/_2774_ ;
wire \myreg/_2775_ ;
wire \myreg/_2776_ ;
wire \myreg/_2777_ ;
wire \myreg/_2778_ ;
wire \myreg/_2779_ ;
wire \myreg/_2780_ ;
wire \myreg/_2781_ ;
wire \myreg/_2782_ ;
wire \myreg/_2783_ ;
wire \myreg/_2784_ ;
wire \myreg/_2785_ ;
wire \myreg/_2786_ ;
wire \myreg/_2787_ ;
wire \myreg/_2788_ ;
wire \myreg/_2789_ ;
wire \myreg/_2790_ ;
wire \myreg/_2791_ ;
wire \myreg/_2792_ ;
wire \myreg/_2793_ ;
wire \myreg/_2794_ ;
wire \myreg/_2795_ ;
wire \myreg/_2796_ ;
wire \myreg/_2797_ ;
wire \myreg/_2798_ ;
wire \myreg/_2799_ ;
wire \myreg/_2800_ ;
wire \myreg/_2801_ ;
wire \myreg/_2802_ ;
wire \myreg/_2803_ ;
wire \myreg/_2804_ ;
wire \myreg/_2805_ ;
wire \myreg/_2806_ ;
wire \myreg/_2807_ ;
wire \myreg/_2808_ ;
wire \myreg/_2809_ ;
wire \myreg/_2810_ ;
wire \myreg/_2811_ ;
wire \myreg/_2812_ ;
wire \myreg/_2813_ ;
wire \myreg/_2814_ ;
wire \myreg/_2815_ ;
wire \myreg/_2816_ ;
wire \myreg/_2817_ ;
wire \myreg/_2818_ ;
wire \myreg/_2819_ ;
wire \myreg/_2820_ ;
wire \myreg/_2821_ ;
wire \myreg/_2822_ ;
wire \myreg/_2823_ ;
wire \myreg/_2824_ ;
wire \myreg/_2825_ ;
wire \myreg/_2826_ ;
wire \myreg/_2827_ ;
wire \myreg/_2828_ ;
wire \myreg/_2829_ ;
wire \myreg/_2830_ ;
wire \myreg/_2831_ ;
wire \myreg/_2832_ ;
wire \myreg/_2833_ ;
wire \myreg/_2834_ ;
wire \myreg/_2835_ ;
wire \myreg/_2836_ ;
wire \myreg/_2837_ ;
wire \myreg/_2838_ ;
wire \myreg/_2839_ ;
wire \myreg/_2840_ ;
wire \myreg/_2841_ ;
wire \myreg/_2842_ ;
wire \myreg/_2843_ ;
wire \myreg/_2844_ ;
wire \myreg/_2845_ ;
wire \myreg/_2846_ ;
wire \myreg/_2847_ ;
wire \myreg/_2848_ ;
wire \myreg/_2849_ ;
wire \myreg/_2850_ ;
wire \myreg/_2851_ ;
wire \myreg/_2852_ ;
wire \myreg/_2853_ ;
wire \myreg/_2854_ ;
wire \myreg/_2855_ ;
wire \myreg/_2856_ ;
wire \myreg/_2857_ ;
wire \myreg/_2858_ ;
wire \myreg/_2859_ ;
wire \myreg/_2860_ ;
wire \myreg/_2861_ ;
wire \myreg/_2862_ ;
wire \myreg/_2863_ ;
wire \myreg/_2864_ ;
wire \myreg/_2865_ ;
wire \myreg/_2866_ ;
wire \myreg/_2867_ ;
wire \myreg/_2868_ ;
wire \myreg/_2869_ ;
wire \myreg/_2870_ ;
wire \myreg/_2871_ ;
wire \myreg/_2872_ ;
wire \myreg/_2873_ ;
wire \myreg/_2874_ ;
wire \myreg/_2875_ ;
wire \myreg/_2876_ ;
wire \myreg/_2877_ ;
wire \myreg/_2878_ ;
wire \myreg/_2879_ ;
wire \myreg/_2880_ ;
wire \myreg/_2881_ ;
wire \myreg/_2882_ ;
wire \myreg/_2883_ ;
wire \myreg/_2884_ ;
wire \myreg/_2885_ ;
wire \myreg/_2886_ ;
wire \myreg/_2887_ ;
wire \myreg/_2888_ ;
wire \myreg/_2889_ ;
wire \myreg/_2890_ ;
wire \myreg/_2891_ ;
wire \myreg/_2892_ ;
wire \myreg/_2893_ ;
wire \myreg/_2894_ ;
wire \myreg/_2895_ ;
wire \myreg/_2896_ ;
wire \myreg/_2897_ ;
wire \myreg/_2898_ ;
wire \myreg/_2899_ ;
wire \myreg/_2900_ ;
wire \myreg/_2901_ ;
wire \myreg/_2902_ ;
wire \myreg/_2903_ ;
wire \myreg/_2904_ ;
wire \myreg/_2905_ ;
wire \myreg/_2906_ ;
wire \myreg/_2907_ ;
wire \myreg/_2908_ ;
wire \myreg/_2909_ ;
wire \myreg/_2910_ ;
wire \myreg/_2911_ ;
wire \myreg/_2912_ ;
wire \myreg/_2913_ ;
wire \myreg/_2914_ ;
wire \myreg/_2915_ ;
wire \myreg/_2916_ ;
wire \myreg/_2917_ ;
wire \myreg/_2918_ ;
wire \myreg/_2919_ ;
wire \myreg/_2920_ ;
wire \myreg/_2921_ ;
wire \myreg/_2922_ ;
wire \myreg/_2923_ ;
wire \myreg/_2924_ ;
wire \myreg/_2925_ ;
wire \myreg/_2926_ ;
wire \myreg/_2927_ ;
wire \myreg/_2928_ ;
wire \myreg/_2929_ ;
wire \myreg/_2930_ ;
wire \myreg/_2931_ ;
wire \myreg/_2932_ ;
wire \myreg/_2933_ ;
wire \myreg/_2934_ ;
wire \myreg/_2935_ ;
wire \myreg/_2936_ ;
wire \myreg/_2937_ ;
wire \myreg/_2938_ ;
wire \myreg/_2939_ ;
wire \myreg/_2940_ ;
wire \myreg/_2941_ ;
wire \myreg/_2942_ ;
wire \myreg/_2943_ ;
wire \myreg/_2944_ ;
wire \myreg/_2945_ ;
wire \myreg/_2946_ ;
wire \myreg/_2947_ ;
wire \myreg/_2948_ ;
wire \myreg/_2949_ ;
wire \myreg/_2950_ ;
wire \myreg/_2951_ ;
wire \myreg/_2952_ ;
wire \myreg/_2953_ ;
wire \myreg/_2954_ ;
wire \myreg/_2955_ ;
wire \myreg/_2956_ ;
wire \myreg/_2957_ ;
wire \myreg/_2958_ ;
wire \myreg/_2959_ ;
wire \myreg/_2960_ ;
wire \myreg/_2961_ ;
wire \myreg/_2962_ ;
wire \myreg/_2963_ ;
wire \myreg/_2964_ ;
wire \myreg/_2965_ ;
wire \myreg/_2966_ ;
wire \myreg/_2967_ ;
wire \myreg/_2968_ ;
wire \myreg/_2969_ ;
wire \myreg/_2970_ ;
wire \myreg/_2971_ ;
wire \myreg/_2972_ ;
wire \myreg/_2973_ ;
wire \myreg/_2974_ ;
wire \myreg/_2975_ ;
wire \myreg/_2976_ ;
wire \myreg/_2977_ ;
wire \myreg/_2978_ ;
wire \myreg/_2979_ ;
wire \myreg/_2980_ ;
wire \myreg/_2981_ ;
wire \myreg/_2982_ ;
wire \myreg/_2983_ ;
wire \myreg/_2984_ ;
wire \myreg/_2985_ ;
wire \myreg/_2986_ ;
wire \myreg/_2987_ ;
wire \myreg/_2988_ ;
wire \myreg/_2989_ ;
wire \myreg/_2990_ ;
wire \myreg/_2991_ ;
wire \myreg/_2992_ ;
wire \myreg/_2993_ ;
wire \myreg/_2994_ ;
wire \myreg/_2995_ ;
wire \myreg/_2996_ ;
wire \myreg/_2997_ ;
wire \myreg/_2998_ ;
wire \myreg/_2999_ ;
wire \myreg/_3000_ ;
wire \myreg/_3001_ ;
wire \myreg/_3002_ ;
wire \myreg/_3003_ ;
wire \myreg/_3004_ ;
wire \myreg/_3005_ ;
wire \myreg/_3006_ ;
wire \myreg/_3007_ ;
wire \myreg/_3008_ ;
wire \myreg/_3009_ ;
wire \myreg/_3010_ ;
wire \myreg/_3011_ ;
wire \myreg/_3012_ ;
wire \myreg/_3013_ ;
wire \myreg/_3014_ ;
wire \myreg/_3015_ ;
wire \myreg/_3016_ ;
wire \myreg/_3017_ ;
wire \myreg/_3018_ ;
wire \myreg/_3019_ ;
wire \myreg/_3020_ ;
wire \myreg/_3021_ ;
wire \myreg/_3022_ ;
wire \myreg/_3023_ ;
wire \myreg/_3024_ ;
wire \myreg/_3025_ ;
wire \myreg/_3026_ ;
wire \myreg/_3027_ ;
wire \myreg/_3028_ ;
wire \myreg/_3029_ ;
wire \myreg/_3030_ ;
wire \myreg/_3031_ ;
wire \myreg/_3032_ ;
wire \myreg/_3033_ ;
wire \myreg/_3034_ ;
wire \myreg/_3035_ ;
wire \myreg/_3036_ ;
wire \myreg/_3037_ ;
wire \myreg/_3038_ ;
wire \myreg/_3039_ ;
wire \myreg/_3040_ ;
wire \myreg/_3041_ ;
wire \myreg/_3042_ ;
wire \myreg/_3043_ ;
wire \myreg/_3044_ ;
wire \myreg/_3045_ ;
wire \myreg/_3046_ ;
wire \myreg/_3047_ ;
wire \myreg/_3048_ ;
wire \myreg/_3049_ ;
wire \myreg/_3050_ ;
wire \myreg/_3051_ ;
wire \myreg/_3052_ ;
wire \myreg/_3053_ ;
wire \myreg/_3054_ ;
wire \myreg/_3055_ ;
wire \myreg/_3056_ ;
wire \myreg/_3057_ ;
wire \myreg/_3058_ ;
wire \myreg/_3059_ ;
wire \myreg/_3060_ ;
wire \myreg/_3061_ ;
wire \myreg/_3062_ ;
wire \myreg/_3063_ ;
wire \myreg/_3064_ ;
wire \myreg/_3065_ ;
wire \myreg/_3066_ ;
wire \myreg/_3067_ ;
wire \myreg/_3068_ ;
wire \myreg/_3069_ ;
wire \myreg/_3070_ ;
wire \myreg/_3071_ ;
wire \myreg/_3072_ ;
wire \myreg/_3073_ ;
wire \myreg/_3074_ ;
wire \myreg/_3075_ ;
wire \myreg/_3076_ ;
wire \myreg/_3077_ ;
wire \myreg/_3078_ ;
wire \myreg/_3079_ ;
wire \myreg/_3080_ ;
wire \myreg/_3081_ ;
wire \myreg/_3082_ ;
wire \myreg/_3083_ ;
wire \myreg/_3084_ ;
wire \myreg/_3085_ ;
wire \myreg/_3086_ ;
wire \myreg/_3087_ ;
wire \myreg/_3088_ ;
wire \myreg/_3089_ ;
wire \myreg/_3090_ ;
wire \myreg/_3091_ ;
wire \myreg/_3092_ ;
wire \myreg/_3093_ ;
wire \myreg/_3094_ ;
wire \myreg/_3095_ ;
wire \myreg/_3096_ ;
wire \myreg/_3097_ ;
wire \myreg/_3098_ ;
wire \myreg/_3099_ ;
wire \myreg/_3100_ ;
wire \myreg/_3101_ ;
wire \myreg/_3102_ ;
wire \myreg/_3103_ ;
wire \myreg/_3104_ ;
wire \myreg/_3105_ ;
wire \myreg/_3106_ ;
wire \myreg/_3107_ ;
wire \myreg/_3108_ ;
wire \myreg/_3109_ ;
wire \myreg/_3110_ ;
wire \myreg/_3111_ ;
wire \myreg/_3112_ ;
wire \myreg/_3113_ ;
wire \myreg/_3114_ ;
wire \myreg/_3115_ ;
wire \myreg/_3116_ ;
wire \myreg/_3117_ ;
wire \myreg/_3118_ ;
wire \myreg/_3119_ ;
wire \myreg/_3120_ ;
wire \myreg/_3121_ ;
wire \myreg/_3122_ ;
wire \myreg/_3123_ ;
wire \myreg/_3124_ ;
wire \myreg/_3125_ ;
wire \myreg/_3126_ ;
wire \myreg/_3127_ ;
wire \myreg/_3128_ ;
wire \myreg/_3129_ ;
wire \myreg/_3130_ ;
wire \myreg/_3131_ ;
wire \myreg/_3132_ ;
wire \myreg/_3133_ ;
wire \myreg/_3134_ ;
wire \myreg/_3135_ ;
wire \myreg/_3136_ ;
wire \myreg/_3137_ ;
wire \myreg/_3138_ ;
wire \myreg/_3139_ ;
wire \myreg/_3140_ ;
wire \myreg/_3141_ ;
wire \myreg/_3142_ ;
wire \myreg/_3143_ ;
wire \myreg/_3144_ ;
wire \myreg/_3145_ ;
wire \myreg/_3146_ ;
wire \myreg/_3147_ ;
wire \myreg/_3148_ ;
wire \myreg/_3149_ ;
wire \myreg/_3150_ ;
wire \myreg/_3151_ ;
wire \myreg/_3152_ ;
wire \myreg/_3153_ ;
wire \myreg/_3154_ ;
wire \myreg/_3155_ ;
wire \myreg/_3156_ ;
wire \myreg/_3157_ ;
wire \myreg/_3158_ ;
wire \myreg/_3159_ ;
wire \myreg/_3160_ ;
wire \myreg/_3161_ ;
wire \myreg/_3162_ ;
wire \myreg/_3163_ ;
wire \myreg/_3164_ ;
wire \myreg/_3165_ ;
wire \myreg/_3166_ ;
wire \myreg/_3167_ ;
wire \myreg/_3168_ ;
wire \myreg/_3169_ ;
wire \myreg/_3170_ ;
wire \myreg/_3171_ ;
wire \myreg/_3172_ ;
wire \myreg/_3173_ ;
wire \myreg/_3174_ ;
wire \myreg/_3175_ ;
wire \myreg/_3176_ ;
wire \myreg/_3177_ ;
wire \myreg/_3178_ ;
wire \myreg/_3179_ ;
wire \myreg/_3180_ ;
wire \myreg/_3181_ ;
wire \myreg/_3182_ ;
wire \myreg/_3183_ ;
wire \myreg/_3184_ ;
wire \myreg/_3185_ ;
wire \myreg/_3186_ ;
wire \myreg/_3187_ ;
wire \myreg/_3188_ ;
wire \myreg/_3189_ ;
wire \myreg/_3190_ ;
wire \myreg/_3191_ ;
wire \myreg/_3192_ ;
wire \myreg/_3193_ ;
wire \myreg/_3194_ ;
wire \myreg/_3195_ ;
wire \myreg/_3196_ ;
wire \myreg/_3197_ ;
wire \myreg/_3198_ ;
wire \myreg/_3199_ ;
wire \myreg/_3200_ ;
wire \myreg/_3201_ ;
wire \myreg/_3202_ ;
wire \myreg/_3203_ ;
wire \myreg/_3204_ ;
wire \myreg/_3205_ ;
wire \myreg/_3206_ ;
wire \myreg/_3207_ ;
wire \myreg/_3208_ ;
wire \myreg/_3209_ ;
wire \myreg/_3210_ ;
wire \myreg/_3211_ ;
wire \myreg/_3212_ ;
wire \myreg/_3213_ ;
wire \myreg/_3214_ ;
wire \myreg/_3215_ ;
wire \myreg/_3216_ ;
wire \myreg/_3217_ ;
wire \myreg/_3218_ ;
wire \myreg/_3219_ ;
wire \myreg/_3220_ ;
wire \myreg/_3221_ ;
wire \myreg/_3222_ ;
wire \myreg/_3223_ ;
wire \myreg/_3224_ ;
wire \myreg/_3225_ ;
wire \myreg/_3226_ ;
wire \myreg/_3227_ ;
wire \myreg/_3228_ ;
wire \myreg/_3229_ ;
wire \myreg/_3230_ ;
wire \myreg/_3231_ ;
wire \myreg/_3232_ ;
wire \myreg/_3233_ ;
wire \myreg/_3234_ ;
wire \myreg/_3235_ ;
wire \myreg/_3236_ ;
wire \myreg/_3237_ ;
wire \myreg/_3238_ ;
wire \myreg/_3239_ ;
wire \myreg/_3240_ ;
wire \myreg/_3241_ ;
wire \myreg/_3242_ ;
wire \myreg/_3243_ ;
wire \myreg/_3244_ ;
wire \myreg/_3245_ ;
wire \myreg/_3246_ ;
wire \myreg/_3247_ ;
wire \myreg/_3248_ ;
wire \myreg/_3249_ ;
wire \myreg/_3250_ ;
wire \myreg/_3251_ ;
wire \myreg/_3252_ ;
wire \myreg/_3253_ ;
wire \myreg/_3254_ ;
wire \myreg/_3255_ ;
wire \myreg/_3256_ ;
wire \myreg/_3257_ ;
wire \myreg/_3258_ ;
wire \myreg/_3259_ ;
wire \myreg/_3260_ ;
wire \myreg/_3261_ ;
wire \myreg/_3262_ ;
wire \myreg/_3263_ ;
wire \myreg/_3264_ ;
wire \myreg/_3265_ ;
wire \myreg/_3266_ ;
wire \myreg/_3267_ ;
wire \myreg/_3268_ ;
wire \myreg/_3269_ ;
wire \myreg/_3270_ ;
wire \myreg/_3271_ ;
wire \myreg/_3272_ ;
wire \myreg/_3273_ ;
wire \myreg/_3274_ ;
wire \myreg/_3275_ ;
wire \myreg/_3276_ ;
wire \myreg/_3277_ ;
wire \myreg/_3278_ ;
wire \myreg/_3279_ ;
wire \myreg/_3280_ ;
wire \myreg/_3281_ ;
wire \myreg/_3282_ ;
wire \myreg/_3283_ ;
wire \myreg/_3284_ ;
wire \myreg/_3285_ ;
wire \myreg/_3286_ ;
wire \myreg/_3287_ ;
wire \myreg/_3288_ ;
wire \myreg/_3289_ ;
wire \myreg/_3290_ ;
wire \myreg/_3291_ ;
wire \myreg/_3292_ ;
wire \myreg/_3293_ ;
wire \myreg/_3294_ ;
wire \myreg/_3295_ ;
wire \myreg/_3296_ ;
wire \myreg/_3297_ ;
wire \myreg/_3298_ ;
wire \myreg/_3299_ ;
wire \myreg/_3300_ ;
wire \myreg/_3301_ ;
wire \myreg/_3302_ ;
wire \myreg/_3303_ ;
wire \myreg/_3304_ ;
wire \myreg/_3305_ ;
wire \myreg/_3306_ ;
wire \myreg/_3307_ ;
wire \myreg/_3308_ ;
wire \myreg/_3309_ ;
wire \myreg/_3310_ ;
wire \myreg/_3311_ ;
wire \myreg/_3312_ ;
wire \myreg/_3313_ ;
wire \myreg/_3314_ ;
wire \myreg/_3315_ ;
wire \myreg/_3316_ ;
wire \myreg/_3317_ ;
wire \myreg/_3318_ ;
wire \myreg/_3319_ ;
wire \myreg/_3320_ ;
wire \myreg/_3321_ ;
wire \myreg/_3322_ ;
wire \myreg/_3323_ ;
wire \myreg/_3324_ ;
wire \myreg/_3325_ ;
wire \myreg/_3326_ ;
wire \myreg/_3327_ ;
wire \myreg/_3328_ ;
wire \myreg/_3329_ ;
wire \myreg/_3330_ ;
wire \myreg/_3331_ ;
wire \myreg/_3332_ ;
wire \myreg/_3333_ ;
wire \myreg/_3334_ ;
wire \myreg/_3335_ ;
wire \myreg/_3336_ ;
wire \myreg/_3337_ ;
wire \myreg/_3338_ ;
wire \myreg/_3339_ ;
wire \myreg/_3340_ ;
wire \myreg/_3341_ ;
wire \myreg/_3342_ ;
wire \myreg/_3343_ ;
wire \myreg/_3344_ ;
wire \myreg/_3345_ ;
wire \myreg/_3346_ ;
wire \myreg/_3347_ ;
wire \myreg/_3348_ ;
wire \myreg/_3349_ ;
wire \myreg/_3350_ ;
wire \myreg/_3351_ ;
wire \myreg/_3352_ ;
wire \myreg/_3353_ ;
wire \myreg/_3354_ ;
wire \myreg/_3355_ ;
wire \myreg/_3356_ ;
wire \myreg/_3357_ ;
wire \myreg/_3358_ ;
wire \myreg/_3359_ ;
wire \myreg/_3360_ ;
wire \myreg/_3361_ ;
wire \myreg/_3362_ ;
wire \myreg/_3363_ ;
wire \myreg/_3364_ ;
wire \myreg/_3365_ ;
wire \myreg/_3366_ ;
wire \myreg/_3367_ ;
wire \myreg/_3368_ ;
wire \myreg/_3369_ ;
wire \myreg/_3370_ ;
wire \myreg/_3371_ ;
wire \myreg/_3372_ ;
wire \myreg/_3373_ ;
wire \myreg/_3374_ ;
wire \myreg/_3375_ ;
wire \myreg/_3376_ ;
wire \myreg/_3377_ ;
wire \myreg/_3378_ ;
wire \myreg/_3379_ ;
wire \myreg/_3380_ ;
wire \myreg/_3381_ ;
wire \myreg/_3382_ ;
wire \myreg/_3383_ ;
wire \myreg/_3384_ ;
wire \myreg/_3385_ ;
wire \myreg/_3386_ ;
wire \myreg/_3387_ ;
wire \myreg/_3388_ ;
wire \myreg/_3389_ ;
wire \myreg/_3390_ ;
wire \myreg/_3391_ ;
wire \myreg/_3392_ ;
wire \myreg/_3393_ ;
wire \myreg/_3394_ ;
wire \myreg/_3395_ ;
wire \myreg/_3396_ ;
wire \myreg/_3397_ ;
wire \myreg/_3398_ ;
wire \myreg/_3399_ ;
wire \myreg/_3400_ ;
wire \myreg/_3401_ ;
wire \myreg/_3402_ ;
wire \myreg/_3403_ ;
wire \myreg/_3404_ ;
wire \myreg/_3405_ ;
wire \myreg/_3406_ ;
wire \myreg/_3407_ ;
wire \myreg/_3408_ ;
wire \myreg/_3409_ ;
wire \myreg/_3410_ ;
wire \myreg/_3411_ ;
wire \myreg/_3412_ ;
wire \myreg/_3413_ ;
wire \myreg/_3414_ ;
wire \myreg/_3415_ ;
wire \myreg/_3416_ ;
wire \myreg/_3417_ ;
wire \myreg/_3418_ ;
wire \myreg/_3419_ ;
wire \myreg/_3420_ ;
wire \myreg/_3421_ ;
wire \myreg/_3422_ ;
wire \myreg/_3423_ ;
wire \myreg/_3424_ ;
wire \myreg/_3425_ ;
wire \myreg/_3426_ ;
wire \myreg/_3427_ ;
wire \myreg/_3428_ ;
wire \myreg/_3429_ ;
wire \myreg/_3430_ ;
wire \myreg/_3431_ ;
wire \myreg/_3432_ ;
wire \myreg/_3433_ ;
wire \myreg/_3434_ ;
wire \myreg/_3435_ ;
wire \myreg/_3436_ ;
wire \myreg/_3437_ ;
wire \myreg/_3438_ ;
wire \myreg/_3439_ ;
wire \myreg/_3440_ ;
wire \myreg/_3441_ ;
wire \myreg/_3442_ ;
wire \myreg/_3443_ ;
wire \myreg/_3444_ ;
wire \myreg/_3445_ ;
wire \myreg/_3446_ ;
wire \myreg/_3447_ ;
wire \myreg/_3448_ ;
wire \myreg/_3449_ ;
wire \myreg/_3450_ ;
wire \myreg/_3451_ ;
wire \myreg/_3452_ ;
wire \myreg/_3453_ ;
wire \myreg/_3454_ ;
wire \myreg/_3455_ ;
wire \myreg/_3456_ ;
wire \myreg/_3457_ ;
wire \myreg/_3458_ ;
wire \myreg/_3459_ ;
wire \myreg/_3460_ ;
wire \myreg/_3461_ ;
wire \myreg/_3462_ ;
wire \myreg/_3463_ ;
wire \myreg/_3464_ ;
wire \myreg/_3465_ ;
wire \myreg/_3466_ ;
wire \myreg/_3467_ ;
wire \myreg/_3468_ ;
wire \myreg/_3469_ ;
wire \myreg/_3470_ ;
wire \myreg/_3471_ ;
wire \myreg/_3472_ ;
wire \myreg/_3473_ ;
wire \myreg/Reg[0][0] ;
wire \myreg/Reg[0][10] ;
wire \myreg/Reg[0][11] ;
wire \myreg/Reg[0][12] ;
wire \myreg/Reg[0][13] ;
wire \myreg/Reg[0][14] ;
wire \myreg/Reg[0][15] ;
wire \myreg/Reg[0][16] ;
wire \myreg/Reg[0][17] ;
wire \myreg/Reg[0][18] ;
wire \myreg/Reg[0][19] ;
wire \myreg/Reg[0][1] ;
wire \myreg/Reg[0][20] ;
wire \myreg/Reg[0][21] ;
wire \myreg/Reg[0][22] ;
wire \myreg/Reg[0][23] ;
wire \myreg/Reg[0][24] ;
wire \myreg/Reg[0][25] ;
wire \myreg/Reg[0][26] ;
wire \myreg/Reg[0][27] ;
wire \myreg/Reg[0][28] ;
wire \myreg/Reg[0][29] ;
wire \myreg/Reg[0][2] ;
wire \myreg/Reg[0][30] ;
wire \myreg/Reg[0][31] ;
wire \myreg/Reg[0][3] ;
wire \myreg/Reg[0][4] ;
wire \myreg/Reg[0][5] ;
wire \myreg/Reg[0][6] ;
wire \myreg/Reg[0][7] ;
wire \myreg/Reg[0][8] ;
wire \myreg/Reg[0][9] ;
wire \myreg/Reg[10][0] ;
wire \myreg/Reg[10][10] ;
wire \myreg/Reg[10][11] ;
wire \myreg/Reg[10][12] ;
wire \myreg/Reg[10][13] ;
wire \myreg/Reg[10][14] ;
wire \myreg/Reg[10][15] ;
wire \myreg/Reg[10][16] ;
wire \myreg/Reg[10][17] ;
wire \myreg/Reg[10][18] ;
wire \myreg/Reg[10][19] ;
wire \myreg/Reg[10][1] ;
wire \myreg/Reg[10][20] ;
wire \myreg/Reg[10][21] ;
wire \myreg/Reg[10][22] ;
wire \myreg/Reg[10][23] ;
wire \myreg/Reg[10][24] ;
wire \myreg/Reg[10][25] ;
wire \myreg/Reg[10][26] ;
wire \myreg/Reg[10][27] ;
wire \myreg/Reg[10][28] ;
wire \myreg/Reg[10][29] ;
wire \myreg/Reg[10][2] ;
wire \myreg/Reg[10][30] ;
wire \myreg/Reg[10][31] ;
wire \myreg/Reg[10][3] ;
wire \myreg/Reg[10][4] ;
wire \myreg/Reg[10][5] ;
wire \myreg/Reg[10][6] ;
wire \myreg/Reg[10][7] ;
wire \myreg/Reg[10][8] ;
wire \myreg/Reg[10][9] ;
wire \myreg/Reg[11][0] ;
wire \myreg/Reg[11][10] ;
wire \myreg/Reg[11][11] ;
wire \myreg/Reg[11][12] ;
wire \myreg/Reg[11][13] ;
wire \myreg/Reg[11][14] ;
wire \myreg/Reg[11][15] ;
wire \myreg/Reg[11][16] ;
wire \myreg/Reg[11][17] ;
wire \myreg/Reg[11][18] ;
wire \myreg/Reg[11][19] ;
wire \myreg/Reg[11][1] ;
wire \myreg/Reg[11][20] ;
wire \myreg/Reg[11][21] ;
wire \myreg/Reg[11][22] ;
wire \myreg/Reg[11][23] ;
wire \myreg/Reg[11][24] ;
wire \myreg/Reg[11][25] ;
wire \myreg/Reg[11][26] ;
wire \myreg/Reg[11][27] ;
wire \myreg/Reg[11][28] ;
wire \myreg/Reg[11][29] ;
wire \myreg/Reg[11][2] ;
wire \myreg/Reg[11][30] ;
wire \myreg/Reg[11][31] ;
wire \myreg/Reg[11][3] ;
wire \myreg/Reg[11][4] ;
wire \myreg/Reg[11][5] ;
wire \myreg/Reg[11][6] ;
wire \myreg/Reg[11][7] ;
wire \myreg/Reg[11][8] ;
wire \myreg/Reg[11][9] ;
wire \myreg/Reg[12][0] ;
wire \myreg/Reg[12][10] ;
wire \myreg/Reg[12][11] ;
wire \myreg/Reg[12][12] ;
wire \myreg/Reg[12][13] ;
wire \myreg/Reg[12][14] ;
wire \myreg/Reg[12][15] ;
wire \myreg/Reg[12][16] ;
wire \myreg/Reg[12][17] ;
wire \myreg/Reg[12][18] ;
wire \myreg/Reg[12][19] ;
wire \myreg/Reg[12][1] ;
wire \myreg/Reg[12][20] ;
wire \myreg/Reg[12][21] ;
wire \myreg/Reg[12][22] ;
wire \myreg/Reg[12][23] ;
wire \myreg/Reg[12][24] ;
wire \myreg/Reg[12][25] ;
wire \myreg/Reg[12][26] ;
wire \myreg/Reg[12][27] ;
wire \myreg/Reg[12][28] ;
wire \myreg/Reg[12][29] ;
wire \myreg/Reg[12][2] ;
wire \myreg/Reg[12][30] ;
wire \myreg/Reg[12][31] ;
wire \myreg/Reg[12][3] ;
wire \myreg/Reg[12][4] ;
wire \myreg/Reg[12][5] ;
wire \myreg/Reg[12][6] ;
wire \myreg/Reg[12][7] ;
wire \myreg/Reg[12][8] ;
wire \myreg/Reg[12][9] ;
wire \myreg/Reg[13][0] ;
wire \myreg/Reg[13][10] ;
wire \myreg/Reg[13][11] ;
wire \myreg/Reg[13][12] ;
wire \myreg/Reg[13][13] ;
wire \myreg/Reg[13][14] ;
wire \myreg/Reg[13][15] ;
wire \myreg/Reg[13][16] ;
wire \myreg/Reg[13][17] ;
wire \myreg/Reg[13][18] ;
wire \myreg/Reg[13][19] ;
wire \myreg/Reg[13][1] ;
wire \myreg/Reg[13][20] ;
wire \myreg/Reg[13][21] ;
wire \myreg/Reg[13][22] ;
wire \myreg/Reg[13][23] ;
wire \myreg/Reg[13][24] ;
wire \myreg/Reg[13][25] ;
wire \myreg/Reg[13][26] ;
wire \myreg/Reg[13][27] ;
wire \myreg/Reg[13][28] ;
wire \myreg/Reg[13][29] ;
wire \myreg/Reg[13][2] ;
wire \myreg/Reg[13][30] ;
wire \myreg/Reg[13][31] ;
wire \myreg/Reg[13][3] ;
wire \myreg/Reg[13][4] ;
wire \myreg/Reg[13][5] ;
wire \myreg/Reg[13][6] ;
wire \myreg/Reg[13][7] ;
wire \myreg/Reg[13][8] ;
wire \myreg/Reg[13][9] ;
wire \myreg/Reg[14][0] ;
wire \myreg/Reg[14][10] ;
wire \myreg/Reg[14][11] ;
wire \myreg/Reg[14][12] ;
wire \myreg/Reg[14][13] ;
wire \myreg/Reg[14][14] ;
wire \myreg/Reg[14][15] ;
wire \myreg/Reg[14][16] ;
wire \myreg/Reg[14][17] ;
wire \myreg/Reg[14][18] ;
wire \myreg/Reg[14][19] ;
wire \myreg/Reg[14][1] ;
wire \myreg/Reg[14][20] ;
wire \myreg/Reg[14][21] ;
wire \myreg/Reg[14][22] ;
wire \myreg/Reg[14][23] ;
wire \myreg/Reg[14][24] ;
wire \myreg/Reg[14][25] ;
wire \myreg/Reg[14][26] ;
wire \myreg/Reg[14][27] ;
wire \myreg/Reg[14][28] ;
wire \myreg/Reg[14][29] ;
wire \myreg/Reg[14][2] ;
wire \myreg/Reg[14][30] ;
wire \myreg/Reg[14][31] ;
wire \myreg/Reg[14][3] ;
wire \myreg/Reg[14][4] ;
wire \myreg/Reg[14][5] ;
wire \myreg/Reg[14][6] ;
wire \myreg/Reg[14][7] ;
wire \myreg/Reg[14][8] ;
wire \myreg/Reg[14][9] ;
wire \myreg/Reg[15][0] ;
wire \myreg/Reg[15][10] ;
wire \myreg/Reg[15][11] ;
wire \myreg/Reg[15][12] ;
wire \myreg/Reg[15][13] ;
wire \myreg/Reg[15][14] ;
wire \myreg/Reg[15][15] ;
wire \myreg/Reg[15][16] ;
wire \myreg/Reg[15][17] ;
wire \myreg/Reg[15][18] ;
wire \myreg/Reg[15][19] ;
wire \myreg/Reg[15][1] ;
wire \myreg/Reg[15][20] ;
wire \myreg/Reg[15][21] ;
wire \myreg/Reg[15][22] ;
wire \myreg/Reg[15][23] ;
wire \myreg/Reg[15][24] ;
wire \myreg/Reg[15][25] ;
wire \myreg/Reg[15][26] ;
wire \myreg/Reg[15][27] ;
wire \myreg/Reg[15][28] ;
wire \myreg/Reg[15][29] ;
wire \myreg/Reg[15][2] ;
wire \myreg/Reg[15][30] ;
wire \myreg/Reg[15][31] ;
wire \myreg/Reg[15][3] ;
wire \myreg/Reg[15][4] ;
wire \myreg/Reg[15][5] ;
wire \myreg/Reg[15][6] ;
wire \myreg/Reg[15][7] ;
wire \myreg/Reg[15][8] ;
wire \myreg/Reg[15][9] ;
wire \myreg/Reg[1][0] ;
wire \myreg/Reg[1][10] ;
wire \myreg/Reg[1][11] ;
wire \myreg/Reg[1][12] ;
wire \myreg/Reg[1][13] ;
wire \myreg/Reg[1][14] ;
wire \myreg/Reg[1][15] ;
wire \myreg/Reg[1][16] ;
wire \myreg/Reg[1][17] ;
wire \myreg/Reg[1][18] ;
wire \myreg/Reg[1][19] ;
wire \myreg/Reg[1][1] ;
wire \myreg/Reg[1][20] ;
wire \myreg/Reg[1][21] ;
wire \myreg/Reg[1][22] ;
wire \myreg/Reg[1][23] ;
wire \myreg/Reg[1][24] ;
wire \myreg/Reg[1][25] ;
wire \myreg/Reg[1][26] ;
wire \myreg/Reg[1][27] ;
wire \myreg/Reg[1][28] ;
wire \myreg/Reg[1][29] ;
wire \myreg/Reg[1][2] ;
wire \myreg/Reg[1][30] ;
wire \myreg/Reg[1][31] ;
wire \myreg/Reg[1][3] ;
wire \myreg/Reg[1][4] ;
wire \myreg/Reg[1][5] ;
wire \myreg/Reg[1][6] ;
wire \myreg/Reg[1][7] ;
wire \myreg/Reg[1][8] ;
wire \myreg/Reg[1][9] ;
wire \myreg/Reg[2][0] ;
wire \myreg/Reg[2][10] ;
wire \myreg/Reg[2][11] ;
wire \myreg/Reg[2][12] ;
wire \myreg/Reg[2][13] ;
wire \myreg/Reg[2][14] ;
wire \myreg/Reg[2][15] ;
wire \myreg/Reg[2][16] ;
wire \myreg/Reg[2][17] ;
wire \myreg/Reg[2][18] ;
wire \myreg/Reg[2][19] ;
wire \myreg/Reg[2][1] ;
wire \myreg/Reg[2][20] ;
wire \myreg/Reg[2][21] ;
wire \myreg/Reg[2][22] ;
wire \myreg/Reg[2][23] ;
wire \myreg/Reg[2][24] ;
wire \myreg/Reg[2][25] ;
wire \myreg/Reg[2][26] ;
wire \myreg/Reg[2][27] ;
wire \myreg/Reg[2][28] ;
wire \myreg/Reg[2][29] ;
wire \myreg/Reg[2][2] ;
wire \myreg/Reg[2][30] ;
wire \myreg/Reg[2][31] ;
wire \myreg/Reg[2][3] ;
wire \myreg/Reg[2][4] ;
wire \myreg/Reg[2][5] ;
wire \myreg/Reg[2][6] ;
wire \myreg/Reg[2][7] ;
wire \myreg/Reg[2][8] ;
wire \myreg/Reg[2][9] ;
wire \myreg/Reg[3][0] ;
wire \myreg/Reg[3][10] ;
wire \myreg/Reg[3][11] ;
wire \myreg/Reg[3][12] ;
wire \myreg/Reg[3][13] ;
wire \myreg/Reg[3][14] ;
wire \myreg/Reg[3][15] ;
wire \myreg/Reg[3][16] ;
wire \myreg/Reg[3][17] ;
wire \myreg/Reg[3][18] ;
wire \myreg/Reg[3][19] ;
wire \myreg/Reg[3][1] ;
wire \myreg/Reg[3][20] ;
wire \myreg/Reg[3][21] ;
wire \myreg/Reg[3][22] ;
wire \myreg/Reg[3][23] ;
wire \myreg/Reg[3][24] ;
wire \myreg/Reg[3][25] ;
wire \myreg/Reg[3][26] ;
wire \myreg/Reg[3][27] ;
wire \myreg/Reg[3][28] ;
wire \myreg/Reg[3][29] ;
wire \myreg/Reg[3][2] ;
wire \myreg/Reg[3][30] ;
wire \myreg/Reg[3][31] ;
wire \myreg/Reg[3][3] ;
wire \myreg/Reg[3][4] ;
wire \myreg/Reg[3][5] ;
wire \myreg/Reg[3][6] ;
wire \myreg/Reg[3][7] ;
wire \myreg/Reg[3][8] ;
wire \myreg/Reg[3][9] ;
wire \myreg/Reg[4][0] ;
wire \myreg/Reg[4][10] ;
wire \myreg/Reg[4][11] ;
wire \myreg/Reg[4][12] ;
wire \myreg/Reg[4][13] ;
wire \myreg/Reg[4][14] ;
wire \myreg/Reg[4][15] ;
wire \myreg/Reg[4][16] ;
wire \myreg/Reg[4][17] ;
wire \myreg/Reg[4][18] ;
wire \myreg/Reg[4][19] ;
wire \myreg/Reg[4][1] ;
wire \myreg/Reg[4][20] ;
wire \myreg/Reg[4][21] ;
wire \myreg/Reg[4][22] ;
wire \myreg/Reg[4][23] ;
wire \myreg/Reg[4][24] ;
wire \myreg/Reg[4][25] ;
wire \myreg/Reg[4][26] ;
wire \myreg/Reg[4][27] ;
wire \myreg/Reg[4][28] ;
wire \myreg/Reg[4][29] ;
wire \myreg/Reg[4][2] ;
wire \myreg/Reg[4][30] ;
wire \myreg/Reg[4][31] ;
wire \myreg/Reg[4][3] ;
wire \myreg/Reg[4][4] ;
wire \myreg/Reg[4][5] ;
wire \myreg/Reg[4][6] ;
wire \myreg/Reg[4][7] ;
wire \myreg/Reg[4][8] ;
wire \myreg/Reg[4][9] ;
wire \myreg/Reg[5][0] ;
wire \myreg/Reg[5][10] ;
wire \myreg/Reg[5][11] ;
wire \myreg/Reg[5][12] ;
wire \myreg/Reg[5][13] ;
wire \myreg/Reg[5][14] ;
wire \myreg/Reg[5][15] ;
wire \myreg/Reg[5][16] ;
wire \myreg/Reg[5][17] ;
wire \myreg/Reg[5][18] ;
wire \myreg/Reg[5][19] ;
wire \myreg/Reg[5][1] ;
wire \myreg/Reg[5][20] ;
wire \myreg/Reg[5][21] ;
wire \myreg/Reg[5][22] ;
wire \myreg/Reg[5][23] ;
wire \myreg/Reg[5][24] ;
wire \myreg/Reg[5][25] ;
wire \myreg/Reg[5][26] ;
wire \myreg/Reg[5][27] ;
wire \myreg/Reg[5][28] ;
wire \myreg/Reg[5][29] ;
wire \myreg/Reg[5][2] ;
wire \myreg/Reg[5][30] ;
wire \myreg/Reg[5][31] ;
wire \myreg/Reg[5][3] ;
wire \myreg/Reg[5][4] ;
wire \myreg/Reg[5][5] ;
wire \myreg/Reg[5][6] ;
wire \myreg/Reg[5][7] ;
wire \myreg/Reg[5][8] ;
wire \myreg/Reg[5][9] ;
wire \myreg/Reg[6][0] ;
wire \myreg/Reg[6][10] ;
wire \myreg/Reg[6][11] ;
wire \myreg/Reg[6][12] ;
wire \myreg/Reg[6][13] ;
wire \myreg/Reg[6][14] ;
wire \myreg/Reg[6][15] ;
wire \myreg/Reg[6][16] ;
wire \myreg/Reg[6][17] ;
wire \myreg/Reg[6][18] ;
wire \myreg/Reg[6][19] ;
wire \myreg/Reg[6][1] ;
wire \myreg/Reg[6][20] ;
wire \myreg/Reg[6][21] ;
wire \myreg/Reg[6][22] ;
wire \myreg/Reg[6][23] ;
wire \myreg/Reg[6][24] ;
wire \myreg/Reg[6][25] ;
wire \myreg/Reg[6][26] ;
wire \myreg/Reg[6][27] ;
wire \myreg/Reg[6][28] ;
wire \myreg/Reg[6][29] ;
wire \myreg/Reg[6][2] ;
wire \myreg/Reg[6][30] ;
wire \myreg/Reg[6][31] ;
wire \myreg/Reg[6][3] ;
wire \myreg/Reg[6][4] ;
wire \myreg/Reg[6][5] ;
wire \myreg/Reg[6][6] ;
wire \myreg/Reg[6][7] ;
wire \myreg/Reg[6][8] ;
wire \myreg/Reg[6][9] ;
wire \myreg/Reg[7][0] ;
wire \myreg/Reg[7][10] ;
wire \myreg/Reg[7][11] ;
wire \myreg/Reg[7][12] ;
wire \myreg/Reg[7][13] ;
wire \myreg/Reg[7][14] ;
wire \myreg/Reg[7][15] ;
wire \myreg/Reg[7][16] ;
wire \myreg/Reg[7][17] ;
wire \myreg/Reg[7][18] ;
wire \myreg/Reg[7][19] ;
wire \myreg/Reg[7][1] ;
wire \myreg/Reg[7][20] ;
wire \myreg/Reg[7][21] ;
wire \myreg/Reg[7][22] ;
wire \myreg/Reg[7][23] ;
wire \myreg/Reg[7][24] ;
wire \myreg/Reg[7][25] ;
wire \myreg/Reg[7][26] ;
wire \myreg/Reg[7][27] ;
wire \myreg/Reg[7][28] ;
wire \myreg/Reg[7][29] ;
wire \myreg/Reg[7][2] ;
wire \myreg/Reg[7][30] ;
wire \myreg/Reg[7][31] ;
wire \myreg/Reg[7][3] ;
wire \myreg/Reg[7][4] ;
wire \myreg/Reg[7][5] ;
wire \myreg/Reg[7][6] ;
wire \myreg/Reg[7][7] ;
wire \myreg/Reg[7][8] ;
wire \myreg/Reg[7][9] ;
wire \myreg/Reg[8][0] ;
wire \myreg/Reg[8][10] ;
wire \myreg/Reg[8][11] ;
wire \myreg/Reg[8][12] ;
wire \myreg/Reg[8][13] ;
wire \myreg/Reg[8][14] ;
wire \myreg/Reg[8][15] ;
wire \myreg/Reg[8][16] ;
wire \myreg/Reg[8][17] ;
wire \myreg/Reg[8][18] ;
wire \myreg/Reg[8][19] ;
wire \myreg/Reg[8][1] ;
wire \myreg/Reg[8][20] ;
wire \myreg/Reg[8][21] ;
wire \myreg/Reg[8][22] ;
wire \myreg/Reg[8][23] ;
wire \myreg/Reg[8][24] ;
wire \myreg/Reg[8][25] ;
wire \myreg/Reg[8][26] ;
wire \myreg/Reg[8][27] ;
wire \myreg/Reg[8][28] ;
wire \myreg/Reg[8][29] ;
wire \myreg/Reg[8][2] ;
wire \myreg/Reg[8][30] ;
wire \myreg/Reg[8][31] ;
wire \myreg/Reg[8][3] ;
wire \myreg/Reg[8][4] ;
wire \myreg/Reg[8][5] ;
wire \myreg/Reg[8][6] ;
wire \myreg/Reg[8][7] ;
wire \myreg/Reg[8][8] ;
wire \myreg/Reg[8][9] ;
wire \myreg/Reg[9][0] ;
wire \myreg/Reg[9][10] ;
wire \myreg/Reg[9][11] ;
wire \myreg/Reg[9][12] ;
wire \myreg/Reg[9][13] ;
wire \myreg/Reg[9][14] ;
wire \myreg/Reg[9][15] ;
wire \myreg/Reg[9][16] ;
wire \myreg/Reg[9][17] ;
wire \myreg/Reg[9][18] ;
wire \myreg/Reg[9][19] ;
wire \myreg/Reg[9][1] ;
wire \myreg/Reg[9][20] ;
wire \myreg/Reg[9][21] ;
wire \myreg/Reg[9][22] ;
wire \myreg/Reg[9][23] ;
wire \myreg/Reg[9][24] ;
wire \myreg/Reg[9][25] ;
wire \myreg/Reg[9][26] ;
wire \myreg/Reg[9][27] ;
wire \myreg/Reg[9][28] ;
wire \myreg/Reg[9][29] ;
wire \myreg/Reg[9][2] ;
wire \myreg/Reg[9][30] ;
wire \myreg/Reg[9][31] ;
wire \myreg/Reg[9][3] ;
wire \myreg/Reg[9][4] ;
wire \myreg/Reg[9][5] ;
wire \myreg/Reg[9][6] ;
wire \myreg/Reg[9][7] ;
wire \myreg/Reg[9][8] ;
wire \myreg/Reg[9][9] ;
wire \mysc/_00_ ;
wire \mysc/_01_ ;
wire \mysc/_02_ ;
wire \mysc/_03_ ;
wire \mysc/_04_ ;
wire \mysc/_05_ ;
wire \mysc/_06_ ;
wire \mysc/_07_ ;
wire \mysc/_08_ ;
wire \mysc/_09_ ;
wire \mysc/_10_ ;
wire \mysc/_11_ ;
wire \mysc/_12_ ;
wire \mysc/_13_ ;
wire \mysc/_14_ ;
wire \mysc/_15_ ;
wire \mysc/_16_ ;
wire \mysc/_17_ ;
wire \mysc/_18_ ;
wire \mysc/_19_ ;
wire \mysc/_20_ ;
wire \mysc/_21_ ;
wire \mysc/_22_ ;
wire \mysc/_23_ ;
wire \mysc/_24_ ;
wire \mysc/_25_ ;
wire \mysc/_26_ ;
wire \mysc/_27_ ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire fanout_net_45 ;
wire fanout_net_46 ;
wire fanout_net_47 ;
wire fanout_net_48 ;
wire fanout_net_49 ;
wire fanout_net_50 ;
wire fanout_net_51 ;
wire fanout_net_52 ;
wire fanout_net_53 ;
wire fanout_net_54 ;
wire fanout_net_55 ;
wire fanout_net_56 ;
wire fanout_net_57 ;
wire fanout_net_58 ;
wire fanout_net_59 ;
wire fanout_net_60 ;
wire fanout_net_61 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [7:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [4:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] araddr_IFU ;
wire [31:0] araddr_LSU ;
wire [31:0] araddr_clint ;
wire [1:0] arburst_IFU ;
wire [1:0] arburst_LSU ;
wire [3:0] arid_IFU ;
wire [3:0] arid_LSU ;
wire [3:0] arid_clint ;
wire [7:0] arlen_IFU ;
wire [7:0] arlen_LSU ;
wire [2:0] arsize_IFU ;
wire [2:0] arsize_LSU ;
wire [31:0] awaddr_LSU ;
wire [1:0] awburst_LSU ;
wire [3:0] awid_LSU ;
wire [7:0] awlen_LSU ;
wire [2:0] awsize_LSU ;
wire [3:0] bid_LSU ;
wire [1:0] bresp_LSU ;
wire [31:0] pc_jump ;
wire [31:0] rdata_IFU ;
wire [31:0] rdata_LSU ;
wire [31:0] rdata_clint ;
wire [3:0] rid_IFU ;
wire [3:0] rid_LSU ;
wire [3:0] rid_clint ;
wire [1:0] rresp_IFU ;
wire [1:0] rresp_LSU ;
wire [1:0] rresp_clint ;
wire [31:0] src1 ;
wire [31:0] src1_raw ;
wire [31:0] src2 ;
wire [31:0] src2_raw ;
wire [31:0] srccs ;
wire [31:0] srccs_raw ;
wire [31:0] wdata_LSU ;
wire [3:0] wstrb_LSU ;
wire [63:0] \myclint/mtime ;
wire [31:0] \myexu/alu_op ;
wire [31:0] \myexu/alu_out ;
wire [2:0] \myidu/state ;
wire [31:0] \myifu/data_out ;
wire [2:0] \myifu/offset ;
wire [2:0] \myifu/state ;
wire [26:0] \myifu/tag_out ;
wire [2:0] \myifu/tmp_offset ;
wire [3:0] \myifu/myicache/valid ;
wire [31:0] \mylsu/araddr_tmp ;
wire [31:0] \mylsu/awaddr_tmp ;
wire [4:0] \mylsu/state ;
wire [2:0] \mylsu/typ_tmp ;
wire [2:0] \myminixbar/state ;
wire [2:0] \mysc/state ;


NAND2_X4 _07_ ( .A1(_03_ ), .A2(_04_ ), .ZN(_05_ ) );
NOR2_X1 _08_ ( .A1(_05_ ), .A2(_02_ ), .ZN(_00_ ) );
XNOR2_X1 _09_ ( .A(_05_ ), .B(_02_ ), .ZN(_01_ ) );
LOGIC0_X1 _10_ ( .Z(_06_ ) );
BUF_X1 _11_ ( .A(fanout_net_1 ), .Z(io_slave_arready ) );
BUF_X1 _12_ ( .A(fanout_net_1 ), .Z(io_slave_awready ) );
BUF_X1 _13_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [0] ) );
BUF_X1 _14_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [1] ) );
BUF_X1 _15_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [2] ) );
BUF_X1 _16_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [3] ) );
BUF_X1 _17_ ( .A(fanout_net_1 ), .Z(\io_slave_bresp [0] ) );
BUF_X1 _18_ ( .A(fanout_net_1 ), .Z(\io_slave_bresp [1] ) );
BUF_X1 _19_ ( .A(fanout_net_1 ), .Z(io_slave_bvalid ) );
BUF_X1 _20_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [0] ) );
BUF_X1 _21_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [1] ) );
BUF_X1 _22_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [2] ) );
BUF_X1 _23_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [3] ) );
BUF_X1 _24_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [4] ) );
BUF_X1 _25_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [5] ) );
BUF_X1 _26_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [6] ) );
BUF_X1 _27_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [7] ) );
BUF_X1 _28_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [8] ) );
BUF_X1 _29_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [9] ) );
BUF_X1 _30_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [10] ) );
BUF_X1 _31_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [11] ) );
BUF_X1 _32_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [12] ) );
BUF_X1 _33_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [13] ) );
BUF_X1 _34_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [14] ) );
BUF_X1 _35_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [15] ) );
BUF_X1 _36_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [16] ) );
BUF_X1 _37_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [17] ) );
BUF_X1 _38_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [18] ) );
BUF_X1 _39_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [19] ) );
BUF_X1 _40_ ( .A(fanout_net_1 ), .Z(\io_slave_rdata [20] ) );
BUF_X1 _41_ ( .A(_06_ ), .Z(\io_slave_rdata [21] ) );
BUF_X1 _42_ ( .A(_06_ ), .Z(\io_slave_rdata [22] ) );
BUF_X1 _43_ ( .A(_06_ ), .Z(\io_slave_rdata [23] ) );
BUF_X1 _44_ ( .A(_06_ ), .Z(\io_slave_rdata [24] ) );
BUF_X1 _45_ ( .A(_06_ ), .Z(\io_slave_rdata [25] ) );
BUF_X1 _46_ ( .A(_06_ ), .Z(\io_slave_rdata [26] ) );
BUF_X1 _47_ ( .A(_06_ ), .Z(\io_slave_rdata [27] ) );
BUF_X1 _48_ ( .A(_06_ ), .Z(\io_slave_rdata [28] ) );
BUF_X1 _49_ ( .A(_06_ ), .Z(\io_slave_rdata [29] ) );
BUF_X1 _50_ ( .A(_06_ ), .Z(\io_slave_rdata [30] ) );
BUF_X1 _51_ ( .A(_06_ ), .Z(\io_slave_rdata [31] ) );
BUF_X1 _52_ ( .A(_06_ ), .Z(\io_slave_rid [0] ) );
BUF_X1 _53_ ( .A(_06_ ), .Z(\io_slave_rid [1] ) );
BUF_X1 _54_ ( .A(_06_ ), .Z(\io_slave_rid [2] ) );
BUF_X1 _55_ ( .A(_06_ ), .Z(\io_slave_rid [3] ) );
BUF_X1 _56_ ( .A(_06_ ), .Z(io_slave_rlast ) );
BUF_X1 _57_ ( .A(_06_ ), .Z(\io_slave_rresp [0] ) );
BUF_X1 _58_ ( .A(_06_ ), .Z(\io_slave_rresp [1] ) );
BUF_X1 _59_ ( .A(_06_ ), .Z(io_slave_rvalid ) );
BUF_X1 _60_ ( .A(_06_ ), .Z(io_slave_wready ) );
BUF_X1 _61_ ( .A(\EX_LS_flag [0] ), .Z(_02_ ) );
BUF_X1 _62_ ( .A(\EX_LS_flag [1] ), .Z(_03_ ) );
BUF_X1 _63_ ( .A(\EX_LS_flag [2] ), .Z(_04_ ) );
BUF_X1 _64_ ( .A(_00_ ), .Z(EX_LS_CSRegWrite ) );
BUF_X1 _65_ ( .A(_01_ ), .Z(EX_LS_RegWrite ) );
MUX2_X1 \myclint/_0526_ ( .A(\myclint/_0068_ ), .B(\myclint/_0093_ ), .S(fanout_net_2 ), .Z(\myclint/_0296_ ) );
MUX2_X1 \myclint/_0527_ ( .A(\myclint/_0079_ ), .B(\myclint/_0094_ ), .S(fanout_net_2 ), .Z(\myclint/_0307_ ) );
MUX2_X1 \myclint/_0528_ ( .A(\myclint/_0090_ ), .B(\myclint/_0095_ ), .S(fanout_net_2 ), .Z(\myclint/_0318_ ) );
MUX2_X1 \myclint/_0529_ ( .A(\myclint/_0101_ ), .B(\myclint/_0096_ ), .S(fanout_net_2 ), .Z(\myclint/_0321_ ) );
MUX2_X1 \myclint/_0530_ ( .A(\myclint/_0112_ ), .B(\myclint/_0097_ ), .S(fanout_net_2 ), .Z(\myclint/_0322_ ) );
MUX2_X1 \myclint/_0531_ ( .A(\myclint/_0123_ ), .B(\myclint/_0098_ ), .S(fanout_net_2 ), .Z(\myclint/_0323_ ) );
MUX2_X1 \myclint/_0532_ ( .A(\myclint/_0128_ ), .B(\myclint/_0099_ ), .S(fanout_net_2 ), .Z(\myclint/_0324_ ) );
MUX2_X1 \myclint/_0533_ ( .A(\myclint/_0129_ ), .B(\myclint/_0100_ ), .S(fanout_net_2 ), .Z(\myclint/_0325_ ) );
MUX2_X1 \myclint/_0534_ ( .A(\myclint/_0130_ ), .B(\myclint/_0102_ ), .S(fanout_net_2 ), .Z(\myclint/_0326_ ) );
MUX2_X1 \myclint/_0535_ ( .A(\myclint/_0131_ ), .B(\myclint/_0103_ ), .S(fanout_net_2 ), .Z(\myclint/_0327_ ) );
MUX2_X1 \myclint/_0536_ ( .A(\myclint/_0069_ ), .B(\myclint/_0104_ ), .S(fanout_net_2 ), .Z(\myclint/_0297_ ) );
MUX2_X1 \myclint/_0537_ ( .A(\myclint/_0070_ ), .B(\myclint/_0105_ ), .S(fanout_net_2 ), .Z(\myclint/_0298_ ) );
MUX2_X1 \myclint/_0538_ ( .A(\myclint/_0071_ ), .B(\myclint/_0106_ ), .S(fanout_net_2 ), .Z(\myclint/_0299_ ) );
MUX2_X1 \myclint/_0539_ ( .A(\myclint/_0072_ ), .B(\myclint/_0107_ ), .S(fanout_net_2 ), .Z(\myclint/_0300_ ) );
MUX2_X1 \myclint/_0540_ ( .A(\myclint/_0073_ ), .B(\myclint/_0108_ ), .S(fanout_net_2 ), .Z(\myclint/_0301_ ) );
MUX2_X1 \myclint/_0541_ ( .A(\myclint/_0074_ ), .B(\myclint/_0109_ ), .S(fanout_net_2 ), .Z(\myclint/_0302_ ) );
MUX2_X1 \myclint/_0542_ ( .A(\myclint/_0075_ ), .B(\myclint/_0110_ ), .S(fanout_net_2 ), .Z(\myclint/_0303_ ) );
MUX2_X1 \myclint/_0543_ ( .A(\myclint/_0076_ ), .B(\myclint/_0111_ ), .S(fanout_net_2 ), .Z(\myclint/_0304_ ) );
MUX2_X1 \myclint/_0544_ ( .A(\myclint/_0077_ ), .B(\myclint/_0113_ ), .S(fanout_net_2 ), .Z(\myclint/_0305_ ) );
MUX2_X1 \myclint/_0545_ ( .A(\myclint/_0078_ ), .B(\myclint/_0114_ ), .S(fanout_net_2 ), .Z(\myclint/_0306_ ) );
MUX2_X1 \myclint/_0546_ ( .A(\myclint/_0080_ ), .B(\myclint/_0115_ ), .S(fanout_net_2 ), .Z(\myclint/_0308_ ) );
MUX2_X1 \myclint/_0547_ ( .A(\myclint/_0081_ ), .B(\myclint/_0116_ ), .S(fanout_net_2 ), .Z(\myclint/_0309_ ) );
MUX2_X1 \myclint/_0548_ ( .A(\myclint/_0082_ ), .B(\myclint/_0117_ ), .S(fanout_net_2 ), .Z(\myclint/_0310_ ) );
MUX2_X1 \myclint/_0549_ ( .A(\myclint/_0083_ ), .B(\myclint/_0118_ ), .S(fanout_net_2 ), .Z(\myclint/_0311_ ) );
MUX2_X1 \myclint/_0550_ ( .A(\myclint/_0084_ ), .B(\myclint/_0119_ ), .S(fanout_net_2 ), .Z(\myclint/_0312_ ) );
MUX2_X1 \myclint/_0551_ ( .A(\myclint/_0085_ ), .B(\myclint/_0120_ ), .S(fanout_net_2 ), .Z(\myclint/_0313_ ) );
MUX2_X1 \myclint/_0552_ ( .A(\myclint/_0086_ ), .B(\myclint/_0121_ ), .S(fanout_net_2 ), .Z(\myclint/_0314_ ) );
MUX2_X1 \myclint/_0553_ ( .A(\myclint/_0087_ ), .B(\myclint/_0122_ ), .S(fanout_net_2 ), .Z(\myclint/_0315_ ) );
MUX2_X1 \myclint/_0554_ ( .A(\myclint/_0088_ ), .B(\myclint/_0124_ ), .S(fanout_net_2 ), .Z(\myclint/_0316_ ) );
MUX2_X1 \myclint/_0555_ ( .A(\myclint/_0089_ ), .B(\myclint/_0125_ ), .S(fanout_net_2 ), .Z(\myclint/_0317_ ) );
MUX2_X1 \myclint/_0556_ ( .A(\myclint/_0091_ ), .B(\myclint/_0126_ ), .S(\myclint/_0000_ ), .Z(\myclint/_0319_ ) );
MUX2_X1 \myclint/_0557_ ( .A(\myclint/_0092_ ), .B(\myclint/_0127_ ), .S(\myclint/_0000_ ), .Z(\myclint/_0320_ ) );
INV_X1 \myclint/_0558_ ( .A(fanout_net_3 ), .ZN(\myclint/_0132_ ) );
BUF_X4 \myclint/_0559_ ( .A(\myclint/_0132_ ), .Z(\myclint/_0133_ ) );
AND2_X1 \myclint/_0560_ ( .A1(\myclint/_0133_ ), .A2(\myclint/_0002_ ), .ZN(\myclint/_0003_ ) );
AND2_X4 \myclint/_0561_ ( .A1(\myclint/_0079_ ), .A2(\myclint/_0068_ ), .ZN(\myclint/_0134_ ) );
NOR2_X1 \myclint/_0562_ ( .A1(\myclint/_0079_ ), .A2(\myclint/_0068_ ), .ZN(\myclint/_0135_ ) );
NOR3_X1 \myclint/_0563_ ( .A1(\myclint/_0134_ ), .A2(\myclint/_0135_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0004_ ) );
AND2_X4 \myclint/_0564_ ( .A1(\myclint/_0134_ ), .A2(\myclint/_0090_ ), .ZN(\myclint/_0136_ ) );
OAI21_X1 \myclint/_0565_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0134_ ), .B2(\myclint/_0090_ ), .ZN(\myclint/_0137_ ) );
NOR2_X1 \myclint/_0566_ ( .A1(\myclint/_0136_ ), .A2(\myclint/_0137_ ), .ZN(\myclint/_0005_ ) );
AND2_X4 \myclint/_0567_ ( .A1(\myclint/_0136_ ), .A2(\myclint/_0101_ ), .ZN(\myclint/_0138_ ) );
AOI21_X1 \myclint/_0568_ ( .A(\myclint/_0101_ ), .B1(\myclint/_0134_ ), .B2(\myclint/_0090_ ), .ZN(\myclint/_0139_ ) );
NOR3_X1 \myclint/_0569_ ( .A1(\myclint/_0138_ ), .A2(fanout_net_3 ), .A3(\myclint/_0139_ ), .ZN(\myclint/_0006_ ) );
AND2_X4 \myclint/_0570_ ( .A1(\myclint/_0138_ ), .A2(\myclint/_0112_ ), .ZN(\myclint/_0140_ ) );
OAI21_X1 \myclint/_0571_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0138_ ), .B2(\myclint/_0112_ ), .ZN(\myclint/_0141_ ) );
NOR2_X1 \myclint/_0572_ ( .A1(\myclint/_0140_ ), .A2(\myclint/_0141_ ), .ZN(\myclint/_0007_ ) );
AND2_X4 \myclint/_0573_ ( .A1(\myclint/_0140_ ), .A2(\myclint/_0123_ ), .ZN(\myclint/_0142_ ) );
AOI21_X1 \myclint/_0574_ ( .A(\myclint/_0123_ ), .B1(\myclint/_0138_ ), .B2(\myclint/_0112_ ), .ZN(\myclint/_0143_ ) );
NOR3_X1 \myclint/_0575_ ( .A1(\myclint/_0142_ ), .A2(fanout_net_3 ), .A3(\myclint/_0143_ ), .ZN(\myclint/_0008_ ) );
AND2_X4 \myclint/_0576_ ( .A1(\myclint/_0142_ ), .A2(\myclint/_0128_ ), .ZN(\myclint/_0144_ ) );
OAI21_X1 \myclint/_0577_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0142_ ), .B2(\myclint/_0128_ ), .ZN(\myclint/_0145_ ) );
NOR2_X1 \myclint/_0578_ ( .A1(\myclint/_0144_ ), .A2(\myclint/_0145_ ), .ZN(\myclint/_0009_ ) );
AND2_X4 \myclint/_0579_ ( .A1(\myclint/_0144_ ), .A2(\myclint/_0129_ ), .ZN(\myclint/_0146_ ) );
AOI21_X1 \myclint/_0580_ ( .A(\myclint/_0129_ ), .B1(\myclint/_0142_ ), .B2(\myclint/_0128_ ), .ZN(\myclint/_0147_ ) );
NOR3_X1 \myclint/_0581_ ( .A1(\myclint/_0146_ ), .A2(fanout_net_3 ), .A3(\myclint/_0147_ ), .ZN(\myclint/_0010_ ) );
AND2_X1 \myclint/_0582_ ( .A1(\myclint/_0146_ ), .A2(\myclint/_0130_ ), .ZN(\myclint/_0148_ ) );
OAI21_X1 \myclint/_0583_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0146_ ), .B2(\myclint/_0130_ ), .ZN(\myclint/_0149_ ) );
NOR2_X1 \myclint/_0584_ ( .A1(\myclint/_0148_ ), .A2(\myclint/_0149_ ), .ZN(\myclint/_0011_ ) );
AND2_X1 \myclint/_0585_ ( .A1(\myclint/_0148_ ), .A2(\myclint/_0131_ ), .ZN(\myclint/_0150_ ) );
AOI21_X1 \myclint/_0586_ ( .A(\myclint/_0131_ ), .B1(\myclint/_0146_ ), .B2(\myclint/_0130_ ), .ZN(\myclint/_0151_ ) );
NOR3_X1 \myclint/_0587_ ( .A1(\myclint/_0150_ ), .A2(fanout_net_3 ), .A3(\myclint/_0151_ ), .ZN(\myclint/_0012_ ) );
AND2_X1 \myclint/_0588_ ( .A1(\myclint/_0150_ ), .A2(\myclint/_0069_ ), .ZN(\myclint/_0152_ ) );
OAI21_X1 \myclint/_0589_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0150_ ), .B2(\myclint/_0069_ ), .ZN(\myclint/_0153_ ) );
NOR2_X1 \myclint/_0590_ ( .A1(\myclint/_0152_ ), .A2(\myclint/_0153_ ), .ZN(\myclint/_0013_ ) );
AOI21_X1 \myclint/_0591_ ( .A(\myclint/_0070_ ), .B1(\myclint/_0150_ ), .B2(\myclint/_0069_ ), .ZN(\myclint/_0154_ ) );
AND2_X1 \myclint/_0592_ ( .A1(\myclint/_0069_ ), .A2(\myclint/_0070_ ), .ZN(\myclint/_0155_ ) );
AND3_X1 \myclint/_0593_ ( .A1(\myclint/_0155_ ), .A2(\myclint/_0130_ ), .A3(\myclint/_0131_ ), .ZN(\myclint/_0156_ ) );
AND2_X1 \myclint/_0594_ ( .A1(\myclint/_0146_ ), .A2(\myclint/_0156_ ), .ZN(\myclint/_0157_ ) );
NOR3_X1 \myclint/_0595_ ( .A1(\myclint/_0154_ ), .A2(fanout_net_3 ), .A3(\myclint/_0157_ ), .ZN(\myclint/_0014_ ) );
AND2_X1 \myclint/_0596_ ( .A1(\myclint/_0157_ ), .A2(\myclint/_0071_ ), .ZN(\myclint/_0158_ ) );
OAI21_X1 \myclint/_0597_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0157_ ), .B2(\myclint/_0071_ ), .ZN(\myclint/_0159_ ) );
NOR2_X1 \myclint/_0598_ ( .A1(\myclint/_0158_ ), .A2(\myclint/_0159_ ), .ZN(\myclint/_0015_ ) );
AND2_X1 \myclint/_0599_ ( .A1(\myclint/_0071_ ), .A2(\myclint/_0072_ ), .ZN(\myclint/_0160_ ) );
AND2_X1 \myclint/_0600_ ( .A1(\myclint/_0157_ ), .A2(\myclint/_0160_ ), .ZN(\myclint/_0161_ ) );
AOI21_X1 \myclint/_0601_ ( .A(\myclint/_0072_ ), .B1(\myclint/_0157_ ), .B2(\myclint/_0071_ ), .ZN(\myclint/_0162_ ) );
NOR3_X1 \myclint/_0602_ ( .A1(\myclint/_0161_ ), .A2(\myclint/_0162_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0016_ ) );
AND2_X1 \myclint/_0603_ ( .A1(\myclint/_0161_ ), .A2(\myclint/_0073_ ), .ZN(\myclint/_0163_ ) );
OAI21_X1 \myclint/_0604_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0161_ ), .B2(\myclint/_0073_ ), .ZN(\myclint/_0164_ ) );
NOR2_X1 \myclint/_0605_ ( .A1(\myclint/_0163_ ), .A2(\myclint/_0164_ ), .ZN(\myclint/_0017_ ) );
AOI21_X1 \myclint/_0606_ ( .A(\myclint/_0074_ ), .B1(\myclint/_0161_ ), .B2(\myclint/_0073_ ), .ZN(\myclint/_0165_ ) );
AND3_X1 \myclint/_0607_ ( .A1(\myclint/_0160_ ), .A2(\myclint/_0073_ ), .A3(\myclint/_0074_ ), .ZN(\myclint/_0166_ ) );
AND4_X1 \myclint/_0608_ ( .A1(\myclint/_0129_ ), .A2(\myclint/_0144_ ), .A3(\myclint/_0156_ ), .A4(\myclint/_0166_ ), .ZN(\myclint/_0167_ ) );
NOR3_X1 \myclint/_0609_ ( .A1(\myclint/_0165_ ), .A2(fanout_net_3 ), .A3(\myclint/_0167_ ), .ZN(\myclint/_0018_ ) );
AND2_X1 \myclint/_0610_ ( .A1(\myclint/_0156_ ), .A2(\myclint/_0166_ ), .ZN(\myclint/_0168_ ) );
AND2_X4 \myclint/_0611_ ( .A1(\myclint/_0146_ ), .A2(\myclint/_0168_ ), .ZN(\myclint/_0169_ ) );
AND2_X1 \myclint/_0612_ ( .A1(\myclint/_0169_ ), .A2(\myclint/_0075_ ), .ZN(\myclint/_0170_ ) );
BUF_X4 \myclint/_0613_ ( .A(\myclint/_0132_ ), .Z(\myclint/_0171_ ) );
OAI21_X1 \myclint/_0614_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0169_ ), .B2(\myclint/_0075_ ), .ZN(\myclint/_0172_ ) );
NOR2_X1 \myclint/_0615_ ( .A1(\myclint/_0170_ ), .A2(\myclint/_0172_ ), .ZN(\myclint/_0019_ ) );
AND2_X1 \myclint/_0616_ ( .A1(\myclint/_0075_ ), .A2(\myclint/_0076_ ), .ZN(\myclint/_0173_ ) );
AND2_X1 \myclint/_0617_ ( .A1(\myclint/_0169_ ), .A2(\myclint/_0173_ ), .ZN(\myclint/_0174_ ) );
AOI21_X1 \myclint/_0618_ ( .A(\myclint/_0076_ ), .B1(\myclint/_0169_ ), .B2(\myclint/_0075_ ), .ZN(\myclint/_0175_ ) );
NOR3_X1 \myclint/_0619_ ( .A1(\myclint/_0174_ ), .A2(\myclint/_0175_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0020_ ) );
AND2_X1 \myclint/_0620_ ( .A1(\myclint/_0174_ ), .A2(\myclint/_0077_ ), .ZN(\myclint/_0176_ ) );
OAI21_X1 \myclint/_0621_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0174_ ), .B2(\myclint/_0077_ ), .ZN(\myclint/_0177_ ) );
NOR2_X1 \myclint/_0622_ ( .A1(\myclint/_0176_ ), .A2(\myclint/_0177_ ), .ZN(\myclint/_0021_ ) );
AOI21_X1 \myclint/_0623_ ( .A(\myclint/_0078_ ), .B1(\myclint/_0174_ ), .B2(\myclint/_0077_ ), .ZN(\myclint/_0178_ ) );
AND3_X1 \myclint/_0624_ ( .A1(\myclint/_0173_ ), .A2(\myclint/_0077_ ), .A3(\myclint/_0078_ ), .ZN(\myclint/_0179_ ) );
AND2_X1 \myclint/_0625_ ( .A1(\myclint/_0169_ ), .A2(\myclint/_0179_ ), .ZN(\myclint/_0180_ ) );
CLKBUF_X2 \myclint/_0626_ ( .A(\myclint/_0180_ ), .Z(\myclint/_0181_ ) );
NOR3_X1 \myclint/_0627_ ( .A1(\myclint/_0178_ ), .A2(fanout_net_3 ), .A3(\myclint/_0181_ ), .ZN(\myclint/_0022_ ) );
AND2_X1 \myclint/_0628_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0080_ ), .ZN(\myclint/_0182_ ) );
OAI21_X1 \myclint/_0629_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0181_ ), .B2(\myclint/_0080_ ), .ZN(\myclint/_0183_ ) );
NOR2_X1 \myclint/_0630_ ( .A1(\myclint/_0182_ ), .A2(\myclint/_0183_ ), .ZN(\myclint/_0023_ ) );
AND2_X1 \myclint/_0631_ ( .A1(\myclint/_0080_ ), .A2(\myclint/_0081_ ), .ZN(\myclint/_0184_ ) );
AND2_X1 \myclint/_0632_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0184_ ), .ZN(\myclint/_0185_ ) );
AOI21_X1 \myclint/_0633_ ( .A(\myclint/_0081_ ), .B1(\myclint/_0181_ ), .B2(\myclint/_0080_ ), .ZN(\myclint/_0186_ ) );
NOR3_X1 \myclint/_0634_ ( .A1(\myclint/_0185_ ), .A2(\myclint/_0186_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0024_ ) );
AND3_X1 \myclint/_0635_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0080_ ), .A3(\myclint/_0081_ ), .ZN(\myclint/_0187_ ) );
AND2_X1 \myclint/_0636_ ( .A1(\myclint/_0187_ ), .A2(\myclint/_0082_ ), .ZN(\myclint/_0188_ ) );
OAI21_X1 \myclint/_0637_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0185_ ), .B2(\myclint/_0082_ ), .ZN(\myclint/_0189_ ) );
NOR2_X1 \myclint/_0638_ ( .A1(\myclint/_0188_ ), .A2(\myclint/_0189_ ), .ZN(\myclint/_0025_ ) );
AOI21_X1 \myclint/_0639_ ( .A(\myclint/_0083_ ), .B1(\myclint/_0185_ ), .B2(\myclint/_0082_ ), .ZN(\myclint/_0190_ ) );
AND3_X1 \myclint/_0640_ ( .A1(\myclint/_0184_ ), .A2(\myclint/_0082_ ), .A3(\myclint/_0083_ ), .ZN(\myclint/_0191_ ) );
AND2_X1 \myclint/_0641_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0191_ ), .ZN(\myclint/_0192_ ) );
NOR3_X1 \myclint/_0642_ ( .A1(\myclint/_0190_ ), .A2(fanout_net_3 ), .A3(\myclint/_0192_ ), .ZN(\myclint/_0026_ ) );
OAI21_X1 \myclint/_0643_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0192_ ), .B2(\myclint/_0084_ ), .ZN(\myclint/_0193_ ) );
AND3_X1 \myclint/_0644_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0084_ ), .A3(\myclint/_0191_ ), .ZN(\myclint/_0194_ ) );
NOR2_X1 \myclint/_0645_ ( .A1(\myclint/_0193_ ), .A2(\myclint/_0194_ ), .ZN(\myclint/_0027_ ) );
AND2_X1 \myclint/_0646_ ( .A1(\myclint/_0179_ ), .A2(\myclint/_0191_ ), .ZN(\myclint/_0195_ ) );
NAND3_X1 \myclint/_0647_ ( .A1(\myclint/_0169_ ), .A2(\myclint/_0084_ ), .A3(\myclint/_0195_ ), .ZN(\myclint/_0196_ ) );
OR2_X1 \myclint/_0648_ ( .A1(\myclint/_0196_ ), .A2(\myclint/_0085_ ), .ZN(\myclint/_0197_ ) );
NAND2_X1 \myclint/_0649_ ( .A1(\myclint/_0196_ ), .A2(\myclint/_0085_ ), .ZN(\myclint/_0198_ ) );
AOI21_X1 \myclint/_0650_ ( .A(fanout_net_3 ), .B1(\myclint/_0197_ ), .B2(\myclint/_0198_ ), .ZN(\myclint/_0028_ ) );
AND2_X1 \myclint/_0651_ ( .A1(\myclint/_0084_ ), .A2(\myclint/_0085_ ), .ZN(\myclint/_0199_ ) );
AND3_X1 \myclint/_0652_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0191_ ), .A3(\myclint/_0199_ ), .ZN(\myclint/_0200_ ) );
AND2_X1 \myclint/_0653_ ( .A1(\myclint/_0200_ ), .A2(\myclint/_0086_ ), .ZN(\myclint/_0201_ ) );
OAI21_X1 \myclint/_0654_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0200_ ), .B2(\myclint/_0086_ ), .ZN(\myclint/_0202_ ) );
NOR2_X1 \myclint/_0655_ ( .A1(\myclint/_0201_ ), .A2(\myclint/_0202_ ), .ZN(\myclint/_0029_ ) );
AOI21_X1 \myclint/_0656_ ( .A(\myclint/_0087_ ), .B1(\myclint/_0200_ ), .B2(\myclint/_0086_ ), .ZN(\myclint/_0203_ ) );
AND2_X1 \myclint/_0657_ ( .A1(\myclint/_0086_ ), .A2(\myclint/_0087_ ), .ZN(\myclint/_0204_ ) );
AND2_X1 \myclint/_0658_ ( .A1(\myclint/_0199_ ), .A2(\myclint/_0204_ ), .ZN(\myclint/_0205_ ) );
AND2_X1 \myclint/_0659_ ( .A1(\myclint/_0191_ ), .A2(\myclint/_0205_ ), .ZN(\myclint/_0206_ ) );
AND2_X1 \myclint/_0660_ ( .A1(\myclint/_0180_ ), .A2(\myclint/_0206_ ), .ZN(\myclint/_0207_ ) );
NOR3_X1 \myclint/_0661_ ( .A1(\myclint/_0203_ ), .A2(fanout_net_3 ), .A3(\myclint/_0207_ ), .ZN(\myclint/_0030_ ) );
OAI21_X1 \myclint/_0662_ ( .A(\myclint/_0133_ ), .B1(\myclint/_0207_ ), .B2(\myclint/_0088_ ), .ZN(\myclint/_0208_ ) );
AND3_X1 \myclint/_0663_ ( .A1(\myclint/_0181_ ), .A2(\myclint/_0088_ ), .A3(\myclint/_0206_ ), .ZN(\myclint/_0209_ ) );
NOR2_X1 \myclint/_0664_ ( .A1(\myclint/_0208_ ), .A2(\myclint/_0209_ ), .ZN(\myclint/_0031_ ) );
AND2_X1 \myclint/_0665_ ( .A1(\myclint/_0088_ ), .A2(\myclint/_0089_ ), .ZN(\myclint/_0210_ ) );
AND2_X1 \myclint/_0666_ ( .A1(\myclint/_0207_ ), .A2(\myclint/_0210_ ), .ZN(\myclint/_0211_ ) );
NOR2_X1 \myclint/_0667_ ( .A1(\myclint/_0209_ ), .A2(\myclint/_0089_ ), .ZN(\myclint/_0212_ ) );
NOR3_X1 \myclint/_0668_ ( .A1(\myclint/_0211_ ), .A2(\myclint/_0212_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0032_ ) );
AND2_X1 \myclint/_0669_ ( .A1(\myclint/_0211_ ), .A2(\myclint/_0091_ ), .ZN(\myclint/_0213_ ) );
OAI21_X1 \myclint/_0670_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0211_ ), .B2(\myclint/_0091_ ), .ZN(\myclint/_0214_ ) );
NOR2_X1 \myclint/_0671_ ( .A1(\myclint/_0213_ ), .A2(\myclint/_0214_ ), .ZN(\myclint/_0033_ ) );
AOI21_X1 \myclint/_0672_ ( .A(\myclint/_0092_ ), .B1(\myclint/_0211_ ), .B2(\myclint/_0091_ ), .ZN(\myclint/_0215_ ) );
AND3_X1 \myclint/_0673_ ( .A1(\myclint/_0210_ ), .A2(\myclint/_0091_ ), .A3(\myclint/_0092_ ), .ZN(\myclint/_0216_ ) );
AND4_X1 \myclint/_0674_ ( .A1(\myclint/_0169_ ), .A2(\myclint/_0179_ ), .A3(\myclint/_0206_ ), .A4(\myclint/_0216_ ), .ZN(\myclint/_0217_ ) );
NOR3_X1 \myclint/_0675_ ( .A1(\myclint/_0215_ ), .A2(fanout_net_3 ), .A3(\myclint/_0217_ ), .ZN(\myclint/_0034_ ) );
AND4_X1 \myclint/_0676_ ( .A1(\myclint/_0179_ ), .A2(\myclint/_0191_ ), .A3(\myclint/_0216_ ), .A4(\myclint/_0205_ ), .ZN(\myclint/_0218_ ) );
AND2_X4 \myclint/_0677_ ( .A1(\myclint/_0169_ ), .A2(\myclint/_0218_ ), .ZN(\myclint/_0219_ ) );
AND2_X4 \myclint/_0678_ ( .A1(\myclint/_0219_ ), .A2(\myclint/_0093_ ), .ZN(\myclint/_0220_ ) );
OAI21_X1 \myclint/_0679_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0219_ ), .B2(\myclint/_0093_ ), .ZN(\myclint/_0221_ ) );
NOR2_X1 \myclint/_0680_ ( .A1(\myclint/_0220_ ), .A2(\myclint/_0221_ ), .ZN(\myclint/_0035_ ) );
AND2_X4 \myclint/_0681_ ( .A1(\myclint/_0220_ ), .A2(\myclint/_0094_ ), .ZN(\myclint/_0222_ ) );
AOI21_X1 \myclint/_0682_ ( .A(\myclint/_0094_ ), .B1(\myclint/_0219_ ), .B2(\myclint/_0093_ ), .ZN(\myclint/_0223_ ) );
NOR3_X1 \myclint/_0683_ ( .A1(\myclint/_0222_ ), .A2(\myclint/_0223_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0036_ ) );
AND2_X4 \myclint/_0684_ ( .A1(\myclint/_0222_ ), .A2(\myclint/_0095_ ), .ZN(\myclint/_0224_ ) );
OAI21_X1 \myclint/_0685_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0222_ ), .B2(\myclint/_0095_ ), .ZN(\myclint/_0225_ ) );
NOR2_X1 \myclint/_0686_ ( .A1(\myclint/_0224_ ), .A2(\myclint/_0225_ ), .ZN(\myclint/_0037_ ) );
AND2_X4 \myclint/_0687_ ( .A1(\myclint/_0224_ ), .A2(\myclint/_0096_ ), .ZN(\myclint/_0226_ ) );
AOI21_X1 \myclint/_0688_ ( .A(\myclint/_0096_ ), .B1(\myclint/_0222_ ), .B2(\myclint/_0095_ ), .ZN(\myclint/_0227_ ) );
NOR3_X1 \myclint/_0689_ ( .A1(\myclint/_0226_ ), .A2(\myclint/_0227_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0038_ ) );
AND2_X4 \myclint/_0690_ ( .A1(\myclint/_0226_ ), .A2(\myclint/_0097_ ), .ZN(\myclint/_0228_ ) );
OAI21_X1 \myclint/_0691_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0226_ ), .B2(\myclint/_0097_ ), .ZN(\myclint/_0229_ ) );
NOR2_X1 \myclint/_0692_ ( .A1(\myclint/_0228_ ), .A2(\myclint/_0229_ ), .ZN(\myclint/_0039_ ) );
AND2_X4 \myclint/_0693_ ( .A1(\myclint/_0228_ ), .A2(\myclint/_0098_ ), .ZN(\myclint/_0230_ ) );
AOI21_X1 \myclint/_0694_ ( .A(\myclint/_0098_ ), .B1(\myclint/_0226_ ), .B2(\myclint/_0097_ ), .ZN(\myclint/_0231_ ) );
NOR3_X1 \myclint/_0695_ ( .A1(\myclint/_0230_ ), .A2(\myclint/_0231_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0040_ ) );
AND2_X4 \myclint/_0696_ ( .A1(\myclint/_0230_ ), .A2(\myclint/_0099_ ), .ZN(\myclint/_0232_ ) );
OAI21_X1 \myclint/_0697_ ( .A(\myclint/_0171_ ), .B1(\myclint/_0230_ ), .B2(\myclint/_0099_ ), .ZN(\myclint/_0233_ ) );
NOR2_X1 \myclint/_0698_ ( .A1(\myclint/_0232_ ), .A2(\myclint/_0233_ ), .ZN(\myclint/_0041_ ) );
AND2_X4 \myclint/_0699_ ( .A1(\myclint/_0232_ ), .A2(\myclint/_0100_ ), .ZN(\myclint/_0234_ ) );
AOI21_X1 \myclint/_0700_ ( .A(\myclint/_0100_ ), .B1(\myclint/_0230_ ), .B2(\myclint/_0099_ ), .ZN(\myclint/_0235_ ) );
NOR3_X1 \myclint/_0701_ ( .A1(\myclint/_0234_ ), .A2(\myclint/_0235_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0042_ ) );
AND2_X1 \myclint/_0702_ ( .A1(\myclint/_0234_ ), .A2(\myclint/_0102_ ), .ZN(\myclint/_0236_ ) );
BUF_X4 \myclint/_0703_ ( .A(\myclint/_0132_ ), .Z(\myclint/_0237_ ) );
OAI21_X1 \myclint/_0704_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0234_ ), .B2(\myclint/_0102_ ), .ZN(\myclint/_0238_ ) );
NOR2_X1 \myclint/_0705_ ( .A1(\myclint/_0236_ ), .A2(\myclint/_0238_ ), .ZN(\myclint/_0043_ ) );
AND2_X1 \myclint/_0706_ ( .A1(\myclint/_0102_ ), .A2(\myclint/_0103_ ), .ZN(\myclint/_0239_ ) );
AND2_X1 \myclint/_0707_ ( .A1(\myclint/_0234_ ), .A2(\myclint/_0239_ ), .ZN(\myclint/_0240_ ) );
AOI21_X1 \myclint/_0708_ ( .A(\myclint/_0103_ ), .B1(\myclint/_0234_ ), .B2(\myclint/_0102_ ), .ZN(\myclint/_0241_ ) );
NOR3_X1 \myclint/_0709_ ( .A1(\myclint/_0240_ ), .A2(\myclint/_0241_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0044_ ) );
AND2_X1 \myclint/_0710_ ( .A1(\myclint/_0240_ ), .A2(\myclint/_0104_ ), .ZN(\myclint/_0242_ ) );
OAI21_X1 \myclint/_0711_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0240_ ), .B2(\myclint/_0104_ ), .ZN(\myclint/_0243_ ) );
NOR2_X1 \myclint/_0712_ ( .A1(\myclint/_0242_ ), .A2(\myclint/_0243_ ), .ZN(\myclint/_0045_ ) );
AOI21_X1 \myclint/_0713_ ( .A(\myclint/_0105_ ), .B1(\myclint/_0240_ ), .B2(\myclint/_0104_ ), .ZN(\myclint/_0244_ ) );
AND3_X1 \myclint/_0714_ ( .A1(\myclint/_0239_ ), .A2(\myclint/_0104_ ), .A3(\myclint/_0105_ ), .ZN(\myclint/_0245_ ) );
AND2_X4 \myclint/_0715_ ( .A1(\myclint/_0234_ ), .A2(\myclint/_0245_ ), .ZN(\myclint/_0246_ ) );
NOR3_X1 \myclint/_0716_ ( .A1(\myclint/_0244_ ), .A2(fanout_net_3 ), .A3(\myclint/_0246_ ), .ZN(\myclint/_0046_ ) );
AND2_X4 \myclint/_0717_ ( .A1(\myclint/_0246_ ), .A2(\myclint/_0106_ ), .ZN(\myclint/_0247_ ) );
OAI21_X1 \myclint/_0718_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0246_ ), .B2(\myclint/_0106_ ), .ZN(\myclint/_0248_ ) );
NOR2_X1 \myclint/_0719_ ( .A1(\myclint/_0247_ ), .A2(\myclint/_0248_ ), .ZN(\myclint/_0047_ ) );
AND2_X4 \myclint/_0720_ ( .A1(\myclint/_0247_ ), .A2(\myclint/_0107_ ), .ZN(\myclint/_0249_ ) );
AOI21_X1 \myclint/_0721_ ( .A(\myclint/_0107_ ), .B1(\myclint/_0246_ ), .B2(\myclint/_0106_ ), .ZN(\myclint/_0250_ ) );
NOR3_X1 \myclint/_0722_ ( .A1(\myclint/_0249_ ), .A2(fanout_net_3 ), .A3(\myclint/_0250_ ), .ZN(\myclint/_0048_ ) );
AND2_X4 \myclint/_0723_ ( .A1(\myclint/_0249_ ), .A2(\myclint/_0108_ ), .ZN(\myclint/_0251_ ) );
OAI21_X1 \myclint/_0724_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0249_ ), .B2(\myclint/_0108_ ), .ZN(\myclint/_0252_ ) );
NOR2_X1 \myclint/_0725_ ( .A1(\myclint/_0251_ ), .A2(\myclint/_0252_ ), .ZN(\myclint/_0049_ ) );
AND2_X4 \myclint/_0726_ ( .A1(\myclint/_0251_ ), .A2(\myclint/_0109_ ), .ZN(\myclint/_0253_ ) );
AOI21_X1 \myclint/_0727_ ( .A(\myclint/_0109_ ), .B1(\myclint/_0249_ ), .B2(\myclint/_0108_ ), .ZN(\myclint/_0254_ ) );
NOR3_X1 \myclint/_0728_ ( .A1(\myclint/_0253_ ), .A2(fanout_net_3 ), .A3(\myclint/_0254_ ), .ZN(\myclint/_0050_ ) );
AND2_X1 \myclint/_0729_ ( .A1(\myclint/_0253_ ), .A2(\myclint/_0110_ ), .ZN(\myclint/_0255_ ) );
OAI21_X1 \myclint/_0730_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0253_ ), .B2(\myclint/_0110_ ), .ZN(\myclint/_0256_ ) );
NOR2_X1 \myclint/_0731_ ( .A1(\myclint/_0255_ ), .A2(\myclint/_0256_ ), .ZN(\myclint/_0051_ ) );
AND2_X1 \myclint/_0732_ ( .A1(\myclint/_0110_ ), .A2(\myclint/_0111_ ), .ZN(\myclint/_0257_ ) );
AND2_X1 \myclint/_0733_ ( .A1(\myclint/_0253_ ), .A2(\myclint/_0257_ ), .ZN(\myclint/_0258_ ) );
AOI21_X1 \myclint/_0734_ ( .A(\myclint/_0111_ ), .B1(\myclint/_0253_ ), .B2(\myclint/_0110_ ), .ZN(\myclint/_0259_ ) );
NOR3_X1 \myclint/_0735_ ( .A1(\myclint/_0258_ ), .A2(\myclint/_0259_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0052_ ) );
AND3_X1 \myclint/_0736_ ( .A1(\myclint/_0253_ ), .A2(\myclint/_0110_ ), .A3(\myclint/_0111_ ), .ZN(\myclint/_0260_ ) );
AND2_X1 \myclint/_0737_ ( .A1(\myclint/_0260_ ), .A2(\myclint/_0113_ ), .ZN(\myclint/_0261_ ) );
OAI21_X1 \myclint/_0738_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0258_ ), .B2(\myclint/_0113_ ), .ZN(\myclint/_0262_ ) );
NOR2_X1 \myclint/_0739_ ( .A1(\myclint/_0261_ ), .A2(\myclint/_0262_ ), .ZN(\myclint/_0053_ ) );
AOI21_X1 \myclint/_0740_ ( .A(\myclint/_0114_ ), .B1(\myclint/_0258_ ), .B2(\myclint/_0113_ ), .ZN(\myclint/_0263_ ) );
AND3_X1 \myclint/_0741_ ( .A1(\myclint/_0257_ ), .A2(\myclint/_0113_ ), .A3(\myclint/_0114_ ), .ZN(\myclint/_0264_ ) );
AND2_X1 \myclint/_0742_ ( .A1(\myclint/_0253_ ), .A2(\myclint/_0264_ ), .ZN(\myclint/_0265_ ) );
NOR3_X1 \myclint/_0743_ ( .A1(\myclint/_0263_ ), .A2(fanout_net_3 ), .A3(\myclint/_0265_ ), .ZN(\myclint/_0054_ ) );
AND2_X1 \myclint/_0744_ ( .A1(\myclint/_0265_ ), .A2(\myclint/_0115_ ), .ZN(\myclint/_0266_ ) );
OAI21_X1 \myclint/_0745_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0265_ ), .B2(\myclint/_0115_ ), .ZN(\myclint/_0267_ ) );
NOR2_X1 \myclint/_0746_ ( .A1(\myclint/_0266_ ), .A2(\myclint/_0267_ ), .ZN(\myclint/_0055_ ) );
AND2_X1 \myclint/_0747_ ( .A1(\myclint/_0115_ ), .A2(\myclint/_0116_ ), .ZN(\myclint/_0268_ ) );
AND2_X1 \myclint/_0748_ ( .A1(\myclint/_0265_ ), .A2(\myclint/_0268_ ), .ZN(\myclint/_0269_ ) );
AOI21_X1 \myclint/_0749_ ( .A(\myclint/_0116_ ), .B1(\myclint/_0265_ ), .B2(\myclint/_0115_ ), .ZN(\myclint/_0270_ ) );
NOR3_X1 \myclint/_0750_ ( .A1(\myclint/_0269_ ), .A2(\myclint/_0270_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0056_ ) );
AND2_X1 \myclint/_0751_ ( .A1(\myclint/_0269_ ), .A2(\myclint/_0117_ ), .ZN(\myclint/_0271_ ) );
OAI21_X1 \myclint/_0752_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0269_ ), .B2(\myclint/_0117_ ), .ZN(\myclint/_0272_ ) );
NOR2_X1 \myclint/_0753_ ( .A1(\myclint/_0271_ ), .A2(\myclint/_0272_ ), .ZN(\myclint/_0057_ ) );
AOI21_X1 \myclint/_0754_ ( .A(\myclint/_0118_ ), .B1(\myclint/_0269_ ), .B2(\myclint/_0117_ ), .ZN(\myclint/_0273_ ) );
AND4_X1 \myclint/_0755_ ( .A1(\myclint/_0117_ ), .A2(\myclint/_0264_ ), .A3(\myclint/_0118_ ), .A4(\myclint/_0268_ ), .ZN(\myclint/_0274_ ) );
AND2_X4 \myclint/_0756_ ( .A1(\myclint/_0253_ ), .A2(\myclint/_0274_ ), .ZN(\myclint/_0275_ ) );
NOR3_X1 \myclint/_0757_ ( .A1(\myclint/_0273_ ), .A2(fanout_net_3 ), .A3(\myclint/_0275_ ), .ZN(\myclint/_0058_ ) );
AND2_X1 \myclint/_0758_ ( .A1(\myclint/_0275_ ), .A2(\myclint/_0119_ ), .ZN(\myclint/_0276_ ) );
OAI21_X1 \myclint/_0759_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0275_ ), .B2(\myclint/_0119_ ), .ZN(\myclint/_0277_ ) );
NOR2_X1 \myclint/_0760_ ( .A1(\myclint/_0276_ ), .A2(\myclint/_0277_ ), .ZN(\myclint/_0059_ ) );
AND2_X4 \myclint/_0761_ ( .A1(\myclint/_0276_ ), .A2(\myclint/_0120_ ), .ZN(\myclint/_0278_ ) );
AOI21_X1 \myclint/_0762_ ( .A(\myclint/_0120_ ), .B1(\myclint/_0275_ ), .B2(\myclint/_0119_ ), .ZN(\myclint/_0279_ ) );
NOR3_X1 \myclint/_0763_ ( .A1(\myclint/_0278_ ), .A2(\myclint/_0279_ ), .A3(fanout_net_3 ), .ZN(\myclint/_0060_ ) );
AND2_X1 \myclint/_0764_ ( .A1(\myclint/_0278_ ), .A2(\myclint/_0121_ ), .ZN(\myclint/_0280_ ) );
OAI21_X1 \myclint/_0765_ ( .A(\myclint/_0237_ ), .B1(\myclint/_0278_ ), .B2(\myclint/_0121_ ), .ZN(\myclint/_0281_ ) );
NOR2_X1 \myclint/_0766_ ( .A1(\myclint/_0280_ ), .A2(\myclint/_0281_ ), .ZN(\myclint/_0061_ ) );
AOI21_X1 \myclint/_0767_ ( .A(\myclint/_0122_ ), .B1(\myclint/_0278_ ), .B2(\myclint/_0121_ ), .ZN(\myclint/_0282_ ) );
AND4_X1 \myclint/_0768_ ( .A1(\myclint/_0120_ ), .A2(\myclint/_0276_ ), .A3(\myclint/_0121_ ), .A4(\myclint/_0122_ ), .ZN(\myclint/_0283_ ) );
NOR3_X1 \myclint/_0769_ ( .A1(\myclint/_0282_ ), .A2(\myclint/_0329_ ), .A3(\myclint/_0283_ ), .ZN(\myclint/_0062_ ) );
AND4_X1 \myclint/_0770_ ( .A1(\myclint/_0119_ ), .A2(\myclint/_0120_ ), .A3(\myclint/_0121_ ), .A4(\myclint/_0122_ ), .ZN(\myclint/_0284_ ) );
AND2_X4 \myclint/_0771_ ( .A1(\myclint/_0275_ ), .A2(\myclint/_0284_ ), .ZN(\myclint/_0285_ ) );
AND2_X1 \myclint/_0772_ ( .A1(\myclint/_0285_ ), .A2(\myclint/_0124_ ), .ZN(\myclint/_0286_ ) );
OAI21_X1 \myclint/_0773_ ( .A(\myclint/_0132_ ), .B1(\myclint/_0285_ ), .B2(\myclint/_0124_ ), .ZN(\myclint/_0287_ ) );
NOR2_X1 \myclint/_0774_ ( .A1(\myclint/_0286_ ), .A2(\myclint/_0287_ ), .ZN(\myclint/_0063_ ) );
AND3_X1 \myclint/_0775_ ( .A1(\myclint/_0285_ ), .A2(\myclint/_0124_ ), .A3(\myclint/_0125_ ), .ZN(\myclint/_0288_ ) );
AOI21_X1 \myclint/_0776_ ( .A(\myclint/_0125_ ), .B1(\myclint/_0285_ ), .B2(\myclint/_0124_ ), .ZN(\myclint/_0289_ ) );
NOR3_X1 \myclint/_0777_ ( .A1(\myclint/_0288_ ), .A2(\myclint/_0289_ ), .A3(\myclint/_0329_ ), .ZN(\myclint/_0064_ ) );
AND3_X4 \myclint/_0778_ ( .A1(\myclint/_0285_ ), .A2(\myclint/_0124_ ), .A3(\myclint/_0125_ ), .ZN(\myclint/_0290_ ) );
AND2_X1 \myclint/_0779_ ( .A1(\myclint/_0290_ ), .A2(\myclint/_0126_ ), .ZN(\myclint/_0291_ ) );
OAI21_X1 \myclint/_0780_ ( .A(\myclint/_0132_ ), .B1(\myclint/_0288_ ), .B2(\myclint/_0126_ ), .ZN(\myclint/_0292_ ) );
NOR2_X1 \myclint/_0781_ ( .A1(\myclint/_0291_ ), .A2(\myclint/_0292_ ), .ZN(\myclint/_0065_ ) );
AND3_X1 \myclint/_0782_ ( .A1(\myclint/_0290_ ), .A2(\myclint/_0126_ ), .A3(\myclint/_0127_ ), .ZN(\myclint/_0293_ ) );
AOI21_X1 \myclint/_0783_ ( .A(\myclint/_0127_ ), .B1(\myclint/_0290_ ), .B2(\myclint/_0126_ ), .ZN(\myclint/_0294_ ) );
NOR3_X1 \myclint/_0784_ ( .A1(\myclint/_0293_ ), .A2(\myclint/_0294_ ), .A3(\myclint/_0329_ ), .ZN(\myclint/_0066_ ) );
NOR2_X1 \myclint/_0785_ ( .A1(\myclint/_0001_ ), .A2(\myclint/_0330_ ), .ZN(\myclint/_0295_ ) );
AOI211_X4 \myclint/_0786_ ( .A(\myclint/_0329_ ), .B(\myclint/_0295_ ), .C1(\myclint/_0328_ ), .C2(\myclint/_0330_ ), .ZN(\myclint/_0067_ ) );
DFF_X1 \myclint/_0787_ ( .D(\myclint/_0461_ ), .CK(clock ), .Q(\myclint/mtime [0] ), .QN(\myclint/_0331_ ) );
DFF_X1 \myclint/_0788_ ( .D(\myclint/_0462_ ), .CK(clock ), .Q(\myclint/mtime [1] ), .QN(\myclint/_0458_ ) );
DFF_X1 \myclint/_0789_ ( .D(\myclint/_0463_ ), .CK(clock ), .Q(\myclint/mtime [2] ), .QN(\myclint/_0457_ ) );
DFF_X1 \myclint/_0790_ ( .D(\myclint/_0464_ ), .CK(clock ), .Q(\myclint/mtime [3] ), .QN(\myclint/_0456_ ) );
DFF_X1 \myclint/_0791_ ( .D(\myclint/_0465_ ), .CK(clock ), .Q(\myclint/mtime [4] ), .QN(\myclint/_0455_ ) );
DFF_X1 \myclint/_0792_ ( .D(\myclint/_0466_ ), .CK(clock ), .Q(\myclint/mtime [5] ), .QN(\myclint/_0454_ ) );
DFF_X1 \myclint/_0793_ ( .D(\myclint/_0467_ ), .CK(clock ), .Q(\myclint/mtime [6] ), .QN(\myclint/_0453_ ) );
DFF_X1 \myclint/_0794_ ( .D(\myclint/_0468_ ), .CK(clock ), .Q(\myclint/mtime [7] ), .QN(\myclint/_0452_ ) );
DFF_X1 \myclint/_0795_ ( .D(\myclint/_0469_ ), .CK(clock ), .Q(\myclint/mtime [8] ), .QN(\myclint/_0451_ ) );
DFF_X1 \myclint/_0796_ ( .D(\myclint/_0470_ ), .CK(clock ), .Q(\myclint/mtime [9] ), .QN(\myclint/_0450_ ) );
DFF_X1 \myclint/_0797_ ( .D(\myclint/_0471_ ), .CK(clock ), .Q(\myclint/mtime [10] ), .QN(\myclint/_0449_ ) );
DFF_X1 \myclint/_0798_ ( .D(\myclint/_0472_ ), .CK(clock ), .Q(\myclint/mtime [11] ), .QN(\myclint/_0448_ ) );
DFF_X1 \myclint/_0799_ ( .D(\myclint/_0473_ ), .CK(clock ), .Q(\myclint/mtime [12] ), .QN(\myclint/_0447_ ) );
DFF_X1 \myclint/_0800_ ( .D(\myclint/_0474_ ), .CK(clock ), .Q(\myclint/mtime [13] ), .QN(\myclint/_0446_ ) );
DFF_X1 \myclint/_0801_ ( .D(\myclint/_0475_ ), .CK(clock ), .Q(\myclint/mtime [14] ), .QN(\myclint/_0445_ ) );
DFF_X1 \myclint/_0802_ ( .D(\myclint/_0476_ ), .CK(clock ), .Q(\myclint/mtime [15] ), .QN(\myclint/_0444_ ) );
DFF_X1 \myclint/_0803_ ( .D(\myclint/_0477_ ), .CK(clock ), .Q(\myclint/mtime [16] ), .QN(\myclint/_0443_ ) );
DFF_X1 \myclint/_0804_ ( .D(\myclint/_0478_ ), .CK(clock ), .Q(\myclint/mtime [17] ), .QN(\myclint/_0442_ ) );
DFF_X1 \myclint/_0805_ ( .D(\myclint/_0479_ ), .CK(clock ), .Q(\myclint/mtime [18] ), .QN(\myclint/_0441_ ) );
DFF_X1 \myclint/_0806_ ( .D(\myclint/_0480_ ), .CK(clock ), .Q(\myclint/mtime [19] ), .QN(\myclint/_0440_ ) );
DFF_X1 \myclint/_0807_ ( .D(\myclint/_0481_ ), .CK(clock ), .Q(\myclint/mtime [20] ), .QN(\myclint/_0439_ ) );
DFF_X1 \myclint/_0808_ ( .D(\myclint/_0482_ ), .CK(clock ), .Q(\myclint/mtime [21] ), .QN(\myclint/_0438_ ) );
DFF_X1 \myclint/_0809_ ( .D(\myclint/_0483_ ), .CK(clock ), .Q(\myclint/mtime [22] ), .QN(\myclint/_0437_ ) );
DFF_X1 \myclint/_0810_ ( .D(\myclint/_0484_ ), .CK(clock ), .Q(\myclint/mtime [23] ), .QN(\myclint/_0436_ ) );
DFF_X1 \myclint/_0811_ ( .D(\myclint/_0485_ ), .CK(clock ), .Q(\myclint/mtime [24] ), .QN(\myclint/_0435_ ) );
DFF_X1 \myclint/_0812_ ( .D(\myclint/_0486_ ), .CK(clock ), .Q(\myclint/mtime [25] ), .QN(\myclint/_0434_ ) );
DFF_X1 \myclint/_0813_ ( .D(\myclint/_0487_ ), .CK(clock ), .Q(\myclint/mtime [26] ), .QN(\myclint/_0433_ ) );
DFF_X1 \myclint/_0814_ ( .D(\myclint/_0488_ ), .CK(clock ), .Q(\myclint/mtime [27] ), .QN(\myclint/_0432_ ) );
DFF_X1 \myclint/_0815_ ( .D(\myclint/_0489_ ), .CK(clock ), .Q(\myclint/mtime [28] ), .QN(\myclint/_0431_ ) );
DFF_X1 \myclint/_0816_ ( .D(\myclint/_0490_ ), .CK(clock ), .Q(\myclint/mtime [29] ), .QN(\myclint/_0430_ ) );
DFF_X1 \myclint/_0817_ ( .D(\myclint/_0491_ ), .CK(clock ), .Q(\myclint/mtime [30] ), .QN(\myclint/_0429_ ) );
DFF_X1 \myclint/_0818_ ( .D(\myclint/_0492_ ), .CK(clock ), .Q(\myclint/mtime [31] ), .QN(\myclint/_0428_ ) );
DFF_X1 \myclint/_0819_ ( .D(\myclint/_0493_ ), .CK(clock ), .Q(\myclint/mtime [32] ), .QN(\myclint/_0427_ ) );
DFF_X1 \myclint/_0820_ ( .D(\myclint/_0494_ ), .CK(clock ), .Q(\myclint/mtime [33] ), .QN(\myclint/_0426_ ) );
DFF_X1 \myclint/_0821_ ( .D(\myclint/_0495_ ), .CK(clock ), .Q(\myclint/mtime [34] ), .QN(\myclint/_0425_ ) );
DFF_X1 \myclint/_0822_ ( .D(\myclint/_0496_ ), .CK(clock ), .Q(\myclint/mtime [35] ), .QN(\myclint/_0424_ ) );
DFF_X1 \myclint/_0823_ ( .D(\myclint/_0497_ ), .CK(clock ), .Q(\myclint/mtime [36] ), .QN(\myclint/_0423_ ) );
DFF_X1 \myclint/_0824_ ( .D(\myclint/_0498_ ), .CK(clock ), .Q(\myclint/mtime [37] ), .QN(\myclint/_0422_ ) );
DFF_X1 \myclint/_0825_ ( .D(\myclint/_0499_ ), .CK(clock ), .Q(\myclint/mtime [38] ), .QN(\myclint/_0421_ ) );
DFF_X1 \myclint/_0826_ ( .D(\myclint/_0500_ ), .CK(clock ), .Q(\myclint/mtime [39] ), .QN(\myclint/_0420_ ) );
DFF_X1 \myclint/_0827_ ( .D(\myclint/_0501_ ), .CK(clock ), .Q(\myclint/mtime [40] ), .QN(\myclint/_0419_ ) );
DFF_X1 \myclint/_0828_ ( .D(\myclint/_0502_ ), .CK(clock ), .Q(\myclint/mtime [41] ), .QN(\myclint/_0418_ ) );
DFF_X1 \myclint/_0829_ ( .D(\myclint/_0503_ ), .CK(clock ), .Q(\myclint/mtime [42] ), .QN(\myclint/_0417_ ) );
DFF_X1 \myclint/_0830_ ( .D(\myclint/_0504_ ), .CK(clock ), .Q(\myclint/mtime [43] ), .QN(\myclint/_0416_ ) );
DFF_X1 \myclint/_0831_ ( .D(\myclint/_0505_ ), .CK(clock ), .Q(\myclint/mtime [44] ), .QN(\myclint/_0415_ ) );
DFF_X1 \myclint/_0832_ ( .D(\myclint/_0506_ ), .CK(clock ), .Q(\myclint/mtime [45] ), .QN(\myclint/_0414_ ) );
DFF_X1 \myclint/_0833_ ( .D(\myclint/_0507_ ), .CK(clock ), .Q(\myclint/mtime [46] ), .QN(\myclint/_0413_ ) );
DFF_X1 \myclint/_0834_ ( .D(\myclint/_0508_ ), .CK(clock ), .Q(\myclint/mtime [47] ), .QN(\myclint/_0412_ ) );
DFF_X1 \myclint/_0835_ ( .D(\myclint/_0509_ ), .CK(clock ), .Q(\myclint/mtime [48] ), .QN(\myclint/_0411_ ) );
DFF_X1 \myclint/_0836_ ( .D(\myclint/_0510_ ), .CK(clock ), .Q(\myclint/mtime [49] ), .QN(\myclint/_0410_ ) );
DFF_X1 \myclint/_0837_ ( .D(\myclint/_0511_ ), .CK(clock ), .Q(\myclint/mtime [50] ), .QN(\myclint/_0409_ ) );
DFF_X1 \myclint/_0838_ ( .D(\myclint/_0512_ ), .CK(clock ), .Q(\myclint/mtime [51] ), .QN(\myclint/_0408_ ) );
DFF_X1 \myclint/_0839_ ( .D(\myclint/_0513_ ), .CK(clock ), .Q(\myclint/mtime [52] ), .QN(\myclint/_0407_ ) );
DFF_X1 \myclint/_0840_ ( .D(\myclint/_0514_ ), .CK(clock ), .Q(\myclint/mtime [53] ), .QN(\myclint/_0406_ ) );
DFF_X1 \myclint/_0841_ ( .D(\myclint/_0515_ ), .CK(clock ), .Q(\myclint/mtime [54] ), .QN(\myclint/_0405_ ) );
DFF_X1 \myclint/_0842_ ( .D(\myclint/_0516_ ), .CK(clock ), .Q(\myclint/mtime [55] ), .QN(\myclint/_0404_ ) );
DFF_X1 \myclint/_0843_ ( .D(\myclint/_0517_ ), .CK(clock ), .Q(\myclint/mtime [56] ), .QN(\myclint/_0403_ ) );
DFF_X1 \myclint/_0844_ ( .D(\myclint/_0518_ ), .CK(clock ), .Q(\myclint/mtime [57] ), .QN(\myclint/_0402_ ) );
DFF_X1 \myclint/_0845_ ( .D(\myclint/_0519_ ), .CK(clock ), .Q(\myclint/mtime [58] ), .QN(\myclint/_0401_ ) );
DFF_X1 \myclint/_0846_ ( .D(\myclint/_0520_ ), .CK(clock ), .Q(\myclint/mtime [59] ), .QN(\myclint/_0400_ ) );
DFF_X1 \myclint/_0847_ ( .D(\myclint/_0521_ ), .CK(clock ), .Q(\myclint/mtime [60] ), .QN(\myclint/_0399_ ) );
DFF_X1 \myclint/_0848_ ( .D(\myclint/_0522_ ), .CK(clock ), .Q(\myclint/mtime [61] ), .QN(\myclint/_0398_ ) );
DFF_X1 \myclint/_0849_ ( .D(\myclint/_0523_ ), .CK(clock ), .Q(\myclint/mtime [62] ), .QN(\myclint/_0397_ ) );
DFF_X1 \myclint/_0850_ ( .D(\myclint/_0524_ ), .CK(clock ), .Q(\myclint/mtime [63] ), .QN(\myclint/_0396_ ) );
DFF_X1 \myclint/_0851_ ( .D(\myclint/_0525_ ), .CK(clock ), .Q(rvalid_clint ), .QN(arready_clint ) );
LOGIC1_X1 \myclint/_0852_ ( .Z(\myclint/_0459_ ) );
LOGIC0_X1 \myclint/_0853_ ( .Z(\myclint/_0460_ ) );
BUF_X1 \myclint/_0854_ ( .A(\myclint/mtime [1] ), .Z(\myclint/_0342_ ) );
BUF_X1 \myclint/_0855_ ( .A(\myclint/mtime [2] ), .Z(\myclint/_0353_ ) );
BUF_X1 \myclint/_0856_ ( .A(\myclint/mtime [3] ), .Z(\myclint/_0364_ ) );
BUF_X1 \myclint/_0857_ ( .A(\myclint/mtime [4] ), .Z(\myclint/_0375_ ) );
BUF_X1 \myclint/_0858_ ( .A(\myclint/mtime [5] ), .Z(\myclint/_0386_ ) );
BUF_X1 \myclint/_0859_ ( .A(\myclint/mtime [6] ), .Z(\myclint/_0391_ ) );
BUF_X1 \myclint/_0860_ ( .A(\myclint/mtime [7] ), .Z(\myclint/_0392_ ) );
BUF_X1 \myclint/_0861_ ( .A(\myclint/mtime [8] ), .Z(\myclint/_0393_ ) );
BUF_X1 \myclint/_0862_ ( .A(\myclint/mtime [9] ), .Z(\myclint/_0394_ ) );
BUF_X1 \myclint/_0863_ ( .A(\myclint/mtime [10] ), .Z(\myclint/_0332_ ) );
BUF_X1 \myclint/_0864_ ( .A(\myclint/mtime [11] ), .Z(\myclint/_0333_ ) );
BUF_X1 \myclint/_0865_ ( .A(\myclint/mtime [12] ), .Z(\myclint/_0334_ ) );
BUF_X1 \myclint/_0866_ ( .A(\myclint/mtime [13] ), .Z(\myclint/_0335_ ) );
BUF_X1 \myclint/_0867_ ( .A(\myclint/mtime [14] ), .Z(\myclint/_0336_ ) );
BUF_X1 \myclint/_0868_ ( .A(\myclint/mtime [15] ), .Z(\myclint/_0337_ ) );
BUF_X1 \myclint/_0869_ ( .A(\myclint/mtime [16] ), .Z(\myclint/_0338_ ) );
BUF_X1 \myclint/_0870_ ( .A(\myclint/mtime [17] ), .Z(\myclint/_0339_ ) );
BUF_X1 \myclint/_0871_ ( .A(\myclint/mtime [18] ), .Z(\myclint/_0340_ ) );
BUF_X1 \myclint/_0872_ ( .A(\myclint/mtime [19] ), .Z(\myclint/_0341_ ) );
BUF_X1 \myclint/_0873_ ( .A(\myclint/mtime [20] ), .Z(\myclint/_0343_ ) );
BUF_X1 \myclint/_0874_ ( .A(\myclint/mtime [21] ), .Z(\myclint/_0344_ ) );
BUF_X1 \myclint/_0875_ ( .A(\myclint/mtime [22] ), .Z(\myclint/_0345_ ) );
BUF_X1 \myclint/_0876_ ( .A(\myclint/mtime [23] ), .Z(\myclint/_0346_ ) );
BUF_X1 \myclint/_0877_ ( .A(\myclint/mtime [24] ), .Z(\myclint/_0347_ ) );
BUF_X1 \myclint/_0878_ ( .A(\myclint/mtime [25] ), .Z(\myclint/_0348_ ) );
BUF_X1 \myclint/_0879_ ( .A(\myclint/mtime [26] ), .Z(\myclint/_0349_ ) );
BUF_X1 \myclint/_0880_ ( .A(\myclint/mtime [27] ), .Z(\myclint/_0350_ ) );
BUF_X1 \myclint/_0881_ ( .A(\myclint/mtime [28] ), .Z(\myclint/_0351_ ) );
BUF_X1 \myclint/_0882_ ( .A(\myclint/mtime [29] ), .Z(\myclint/_0352_ ) );
BUF_X1 \myclint/_0883_ ( .A(\myclint/mtime [30] ), .Z(\myclint/_0354_ ) );
BUF_X1 \myclint/_0884_ ( .A(\myclint/mtime [31] ), .Z(\myclint/_0355_ ) );
BUF_X1 \myclint/_0885_ ( .A(\myclint/mtime [32] ), .Z(\myclint/_0356_ ) );
BUF_X1 \myclint/_0886_ ( .A(\myclint/mtime [33] ), .Z(\myclint/_0357_ ) );
BUF_X1 \myclint/_0887_ ( .A(\myclint/mtime [34] ), .Z(\myclint/_0358_ ) );
BUF_X1 \myclint/_0888_ ( .A(\myclint/mtime [35] ), .Z(\myclint/_0359_ ) );
BUF_X1 \myclint/_0889_ ( .A(\myclint/mtime [36] ), .Z(\myclint/_0360_ ) );
BUF_X1 \myclint/_0890_ ( .A(\myclint/mtime [37] ), .Z(\myclint/_0361_ ) );
BUF_X1 \myclint/_0891_ ( .A(\myclint/mtime [38] ), .Z(\myclint/_0362_ ) );
BUF_X1 \myclint/_0892_ ( .A(\myclint/mtime [39] ), .Z(\myclint/_0363_ ) );
BUF_X1 \myclint/_0893_ ( .A(\myclint/mtime [40] ), .Z(\myclint/_0365_ ) );
BUF_X1 \myclint/_0894_ ( .A(\myclint/mtime [41] ), .Z(\myclint/_0366_ ) );
BUF_X1 \myclint/_0895_ ( .A(\myclint/mtime [42] ), .Z(\myclint/_0367_ ) );
BUF_X1 \myclint/_0896_ ( .A(\myclint/mtime [43] ), .Z(\myclint/_0368_ ) );
BUF_X1 \myclint/_0897_ ( .A(\myclint/mtime [44] ), .Z(\myclint/_0369_ ) );
BUF_X1 \myclint/_0898_ ( .A(\myclint/mtime [45] ), .Z(\myclint/_0370_ ) );
BUF_X1 \myclint/_0899_ ( .A(\myclint/mtime [46] ), .Z(\myclint/_0371_ ) );
BUF_X1 \myclint/_0900_ ( .A(\myclint/mtime [47] ), .Z(\myclint/_0372_ ) );
BUF_X1 \myclint/_0901_ ( .A(\myclint/mtime [48] ), .Z(\myclint/_0373_ ) );
BUF_X1 \myclint/_0902_ ( .A(\myclint/mtime [49] ), .Z(\myclint/_0374_ ) );
BUF_X1 \myclint/_0903_ ( .A(\myclint/mtime [50] ), .Z(\myclint/_0376_ ) );
BUF_X1 \myclint/_0904_ ( .A(\myclint/mtime [51] ), .Z(\myclint/_0377_ ) );
BUF_X1 \myclint/_0905_ ( .A(\myclint/mtime [52] ), .Z(\myclint/_0378_ ) );
BUF_X1 \myclint/_0906_ ( .A(\myclint/mtime [53] ), .Z(\myclint/_0379_ ) );
BUF_X1 \myclint/_0907_ ( .A(\myclint/mtime [54] ), .Z(\myclint/_0380_ ) );
BUF_X1 \myclint/_0908_ ( .A(\myclint/mtime [55] ), .Z(\myclint/_0381_ ) );
BUF_X1 \myclint/_0909_ ( .A(\myclint/mtime [56] ), .Z(\myclint/_0382_ ) );
BUF_X1 \myclint/_0910_ ( .A(\myclint/mtime [57] ), .Z(\myclint/_0383_ ) );
BUF_X1 \myclint/_0911_ ( .A(\myclint/mtime [58] ), .Z(\myclint/_0384_ ) );
BUF_X1 \myclint/_0912_ ( .A(\myclint/mtime [59] ), .Z(\myclint/_0385_ ) );
BUF_X1 \myclint/_0913_ ( .A(\myclint/mtime [60] ), .Z(\myclint/_0387_ ) );
BUF_X1 \myclint/_0914_ ( .A(\myclint/mtime [61] ), .Z(\myclint/_0388_ ) );
BUF_X1 \myclint/_0915_ ( .A(\myclint/mtime [62] ), .Z(\myclint/_0389_ ) );
BUF_X1 \myclint/_0916_ ( .A(\myclint/mtime [63] ), .Z(\myclint/_0390_ ) );
BUF_X1 \myclint/_0917_ ( .A(\myclint/_0331_ ), .Z(\myclint/_0395_ ) );
BUF_X1 \myclint/_0918_ ( .A(\arid_clint [0] ), .Z(\rid_clint [0] ) );
BUF_X1 \myclint/_0919_ ( .A(\arid_clint [1] ), .Z(\rid_clint [1] ) );
BUF_X1 \myclint/_0920_ ( .A(\arid_clint [2] ), .Z(\rid_clint [2] ) );
BUF_X1 \myclint/_0921_ ( .A(\arid_clint [3] ), .Z(\rid_clint [3] ) );
BUF_X1 \myclint/_0922_ ( .A(\myclint/_0459_ ), .Z(rlast_clint ) );
BUF_X1 \myclint/_0923_ ( .A(\myclint/_0460_ ), .Z(\rresp_clint [0] ) );
BUF_X1 \myclint/_0924_ ( .A(\myclint/_0460_ ), .Z(\rresp_clint [1] ) );
BUF_X1 \myclint/_0925_ ( .A(\myclint/mtime [1] ), .Z(\myclint/_0079_ ) );
BUF_X1 \myclint/_0926_ ( .A(\myclint/mtime [0] ), .Z(\myclint/_0068_ ) );
BUF_X1 \myclint/_0927_ ( .A(\myclint/mtime [2] ), .Z(\myclint/_0090_ ) );
BUF_X1 \myclint/_0928_ ( .A(\myclint/mtime [3] ), .Z(\myclint/_0101_ ) );
BUF_X1 \myclint/_0929_ ( .A(\myclint/mtime [4] ), .Z(\myclint/_0112_ ) );
BUF_X1 \myclint/_0930_ ( .A(\myclint/mtime [5] ), .Z(\myclint/_0123_ ) );
BUF_X1 \myclint/_0931_ ( .A(\myclint/mtime [6] ), .Z(\myclint/_0128_ ) );
BUF_X1 \myclint/_0932_ ( .A(\myclint/mtime [7] ), .Z(\myclint/_0129_ ) );
BUF_X1 \myclint/_0933_ ( .A(\myclint/mtime [8] ), .Z(\myclint/_0130_ ) );
BUF_X1 \myclint/_0934_ ( .A(\myclint/mtime [9] ), .Z(\myclint/_0131_ ) );
BUF_X1 \myclint/_0935_ ( .A(\myclint/mtime [10] ), .Z(\myclint/_0069_ ) );
BUF_X1 \myclint/_0936_ ( .A(\myclint/mtime [11] ), .Z(\myclint/_0070_ ) );
BUF_X1 \myclint/_0937_ ( .A(\myclint/mtime [12] ), .Z(\myclint/_0071_ ) );
BUF_X1 \myclint/_0938_ ( .A(\myclint/mtime [13] ), .Z(\myclint/_0072_ ) );
BUF_X1 \myclint/_0939_ ( .A(\myclint/mtime [14] ), .Z(\myclint/_0073_ ) );
BUF_X1 \myclint/_0940_ ( .A(\myclint/mtime [15] ), .Z(\myclint/_0074_ ) );
BUF_X1 \myclint/_0941_ ( .A(\myclint/mtime [16] ), .Z(\myclint/_0075_ ) );
BUF_X1 \myclint/_0942_ ( .A(\myclint/mtime [17] ), .Z(\myclint/_0076_ ) );
BUF_X1 \myclint/_0943_ ( .A(\myclint/mtime [18] ), .Z(\myclint/_0077_ ) );
BUF_X1 \myclint/_0944_ ( .A(\myclint/mtime [19] ), .Z(\myclint/_0078_ ) );
BUF_X1 \myclint/_0945_ ( .A(\myclint/mtime [20] ), .Z(\myclint/_0080_ ) );
BUF_X1 \myclint/_0946_ ( .A(\myclint/mtime [21] ), .Z(\myclint/_0081_ ) );
BUF_X1 \myclint/_0947_ ( .A(\myclint/mtime [22] ), .Z(\myclint/_0082_ ) );
BUF_X1 \myclint/_0948_ ( .A(\myclint/mtime [23] ), .Z(\myclint/_0083_ ) );
BUF_X1 \myclint/_0949_ ( .A(\myclint/mtime [24] ), .Z(\myclint/_0084_ ) );
BUF_X1 \myclint/_0950_ ( .A(\myclint/mtime [25] ), .Z(\myclint/_0085_ ) );
BUF_X1 \myclint/_0951_ ( .A(\myclint/mtime [26] ), .Z(\myclint/_0086_ ) );
BUF_X1 \myclint/_0952_ ( .A(\myclint/mtime [27] ), .Z(\myclint/_0087_ ) );
BUF_X1 \myclint/_0953_ ( .A(\myclint/mtime [28] ), .Z(\myclint/_0088_ ) );
BUF_X1 \myclint/_0954_ ( .A(\myclint/mtime [29] ), .Z(\myclint/_0089_ ) );
BUF_X1 \myclint/_0955_ ( .A(\myclint/mtime [30] ), .Z(\myclint/_0091_ ) );
BUF_X1 \myclint/_0956_ ( .A(\myclint/mtime [31] ), .Z(\myclint/_0092_ ) );
BUF_X1 \myclint/_0957_ ( .A(\myclint/mtime [32] ), .Z(\myclint/_0093_ ) );
BUF_X1 \myclint/_0958_ ( .A(\myclint/mtime [33] ), .Z(\myclint/_0094_ ) );
BUF_X1 \myclint/_0959_ ( .A(\myclint/mtime [34] ), .Z(\myclint/_0095_ ) );
BUF_X1 \myclint/_0960_ ( .A(\myclint/mtime [35] ), .Z(\myclint/_0096_ ) );
BUF_X1 \myclint/_0961_ ( .A(\myclint/mtime [36] ), .Z(\myclint/_0097_ ) );
BUF_X1 \myclint/_0962_ ( .A(\myclint/mtime [37] ), .Z(\myclint/_0098_ ) );
BUF_X1 \myclint/_0963_ ( .A(\myclint/mtime [38] ), .Z(\myclint/_0099_ ) );
BUF_X1 \myclint/_0964_ ( .A(\myclint/mtime [39] ), .Z(\myclint/_0100_ ) );
BUF_X1 \myclint/_0965_ ( .A(\myclint/mtime [40] ), .Z(\myclint/_0102_ ) );
BUF_X1 \myclint/_0966_ ( .A(\myclint/mtime [41] ), .Z(\myclint/_0103_ ) );
BUF_X1 \myclint/_0967_ ( .A(\myclint/mtime [42] ), .Z(\myclint/_0104_ ) );
BUF_X1 \myclint/_0968_ ( .A(\myclint/mtime [43] ), .Z(\myclint/_0105_ ) );
BUF_X1 \myclint/_0969_ ( .A(\myclint/mtime [44] ), .Z(\myclint/_0106_ ) );
BUF_X1 \myclint/_0970_ ( .A(\myclint/mtime [45] ), .Z(\myclint/_0107_ ) );
BUF_X1 \myclint/_0971_ ( .A(\myclint/mtime [46] ), .Z(\myclint/_0108_ ) );
BUF_X1 \myclint/_0972_ ( .A(\myclint/mtime [47] ), .Z(\myclint/_0109_ ) );
BUF_X1 \myclint/_0973_ ( .A(\myclint/mtime [48] ), .Z(\myclint/_0110_ ) );
BUF_X1 \myclint/_0974_ ( .A(\myclint/mtime [49] ), .Z(\myclint/_0111_ ) );
BUF_X1 \myclint/_0975_ ( .A(\myclint/mtime [50] ), .Z(\myclint/_0113_ ) );
BUF_X1 \myclint/_0976_ ( .A(\myclint/mtime [51] ), .Z(\myclint/_0114_ ) );
BUF_X1 \myclint/_0977_ ( .A(\myclint/mtime [52] ), .Z(\myclint/_0115_ ) );
BUF_X1 \myclint/_0978_ ( .A(\myclint/mtime [53] ), .Z(\myclint/_0116_ ) );
BUF_X1 \myclint/_0979_ ( .A(\myclint/mtime [54] ), .Z(\myclint/_0117_ ) );
BUF_X1 \myclint/_0980_ ( .A(\myclint/mtime [55] ), .Z(\myclint/_0118_ ) );
BUF_X1 \myclint/_0981_ ( .A(\myclint/mtime [56] ), .Z(\myclint/_0119_ ) );
BUF_X1 \myclint/_0982_ ( .A(\myclint/mtime [57] ), .Z(\myclint/_0120_ ) );
BUF_X1 \myclint/_0983_ ( .A(\myclint/mtime [58] ), .Z(\myclint/_0121_ ) );
BUF_X1 \myclint/_0984_ ( .A(\myclint/mtime [59] ), .Z(\myclint/_0122_ ) );
BUF_X1 \myclint/_0985_ ( .A(\myclint/mtime [60] ), .Z(\myclint/_0124_ ) );
BUF_X1 \myclint/_0986_ ( .A(\myclint/mtime [61] ), .Z(\myclint/_0125_ ) );
BUF_X1 \myclint/_0987_ ( .A(\myclint/mtime [62] ), .Z(\myclint/_0126_ ) );
BUF_X1 \myclint/_0988_ ( .A(\myclint/mtime [63] ), .Z(\myclint/_0127_ ) );
BUF_X1 \myclint/_0989_ ( .A(rready_clint ), .Z(\myclint/_0328_ ) );
BUF_X1 \myclint/_0990_ ( .A(arvalid_clint ), .Z(\myclint/_0001_ ) );
BUF_X1 \myclint/_0991_ ( .A(rvalid_clint ), .Z(\myclint/_0330_ ) );
BUF_X1 \myclint/_0992_ ( .A(\araddr_clint [2] ), .Z(\myclint/_0000_ ) );
BUF_X1 \myclint/_0993_ ( .A(\myclint/_0296_ ), .Z(\rdata_clint [0] ) );
BUF_X1 \myclint/_0994_ ( .A(\myclint/_0307_ ), .Z(\rdata_clint [1] ) );
BUF_X1 \myclint/_0995_ ( .A(\myclint/_0318_ ), .Z(\rdata_clint [2] ) );
BUF_X1 \myclint/_0996_ ( .A(\myclint/_0321_ ), .Z(\rdata_clint [3] ) );
BUF_X1 \myclint/_0997_ ( .A(\myclint/_0322_ ), .Z(\rdata_clint [4] ) );
BUF_X1 \myclint/_0998_ ( .A(\myclint/_0323_ ), .Z(\rdata_clint [5] ) );
BUF_X1 \myclint/_0999_ ( .A(\myclint/_0324_ ), .Z(\rdata_clint [6] ) );
BUF_X1 \myclint/_1000_ ( .A(\myclint/_0325_ ), .Z(\rdata_clint [7] ) );
BUF_X1 \myclint/_1001_ ( .A(\myclint/_0326_ ), .Z(\rdata_clint [8] ) );
BUF_X1 \myclint/_1002_ ( .A(\myclint/_0327_ ), .Z(\rdata_clint [9] ) );
BUF_X1 \myclint/_1003_ ( .A(\myclint/_0297_ ), .Z(\rdata_clint [10] ) );
BUF_X1 \myclint/_1004_ ( .A(\myclint/_0298_ ), .Z(\rdata_clint [11] ) );
BUF_X1 \myclint/_1005_ ( .A(\myclint/_0299_ ), .Z(\rdata_clint [12] ) );
BUF_X1 \myclint/_1006_ ( .A(\myclint/_0300_ ), .Z(\rdata_clint [13] ) );
BUF_X1 \myclint/_1007_ ( .A(\myclint/_0301_ ), .Z(\rdata_clint [14] ) );
BUF_X1 \myclint/_1008_ ( .A(\myclint/_0302_ ), .Z(\rdata_clint [15] ) );
BUF_X1 \myclint/_1009_ ( .A(\myclint/_0303_ ), .Z(\rdata_clint [16] ) );
BUF_X1 \myclint/_1010_ ( .A(\myclint/_0304_ ), .Z(\rdata_clint [17] ) );
BUF_X1 \myclint/_1011_ ( .A(\myclint/_0305_ ), .Z(\rdata_clint [18] ) );
BUF_X1 \myclint/_1012_ ( .A(\myclint/_0306_ ), .Z(\rdata_clint [19] ) );
BUF_X1 \myclint/_1013_ ( .A(\myclint/_0308_ ), .Z(\rdata_clint [20] ) );
BUF_X1 \myclint/_1014_ ( .A(\myclint/_0309_ ), .Z(\rdata_clint [21] ) );
BUF_X1 \myclint/_1015_ ( .A(\myclint/_0310_ ), .Z(\rdata_clint [22] ) );
BUF_X1 \myclint/_1016_ ( .A(\myclint/_0311_ ), .Z(\rdata_clint [23] ) );
BUF_X1 \myclint/_1017_ ( .A(\myclint/_0312_ ), .Z(\rdata_clint [24] ) );
BUF_X1 \myclint/_1018_ ( .A(\myclint/_0313_ ), .Z(\rdata_clint [25] ) );
BUF_X1 \myclint/_1019_ ( .A(\myclint/_0314_ ), .Z(\rdata_clint [26] ) );
BUF_X1 \myclint/_1020_ ( .A(\myclint/_0315_ ), .Z(\rdata_clint [27] ) );
BUF_X1 \myclint/_1021_ ( .A(\myclint/_0316_ ), .Z(\rdata_clint [28] ) );
BUF_X1 \myclint/_1022_ ( .A(\myclint/_0317_ ), .Z(\rdata_clint [29] ) );
BUF_X1 \myclint/_1023_ ( .A(\myclint/_0319_ ), .Z(\rdata_clint [30] ) );
BUF_X1 \myclint/_1024_ ( .A(\myclint/_0320_ ), .Z(\rdata_clint [31] ) );
BUF_X1 \myclint/_1025_ ( .A(\myclint/_0331_ ), .Z(\myclint/_0002_ ) );
BUF_X1 \myclint/_1026_ ( .A(reset ), .Z(\myclint/_0329_ ) );
BUF_X1 \myclint/_1027_ ( .A(\myclint/_0003_ ), .Z(\myclint/_0461_ ) );
BUF_X1 \myclint/_1028_ ( .A(\myclint/_0004_ ), .Z(\myclint/_0462_ ) );
BUF_X1 \myclint/_1029_ ( .A(\myclint/_0005_ ), .Z(\myclint/_0463_ ) );
BUF_X1 \myclint/_1030_ ( .A(\myclint/_0006_ ), .Z(\myclint/_0464_ ) );
BUF_X1 \myclint/_1031_ ( .A(\myclint/_0007_ ), .Z(\myclint/_0465_ ) );
BUF_X1 \myclint/_1032_ ( .A(\myclint/_0008_ ), .Z(\myclint/_0466_ ) );
BUF_X1 \myclint/_1033_ ( .A(\myclint/_0009_ ), .Z(\myclint/_0467_ ) );
BUF_X1 \myclint/_1034_ ( .A(\myclint/_0010_ ), .Z(\myclint/_0468_ ) );
BUF_X1 \myclint/_1035_ ( .A(\myclint/_0011_ ), .Z(\myclint/_0469_ ) );
BUF_X1 \myclint/_1036_ ( .A(\myclint/_0012_ ), .Z(\myclint/_0470_ ) );
BUF_X1 \myclint/_1037_ ( .A(\myclint/_0013_ ), .Z(\myclint/_0471_ ) );
BUF_X1 \myclint/_1038_ ( .A(\myclint/_0014_ ), .Z(\myclint/_0472_ ) );
BUF_X1 \myclint/_1039_ ( .A(\myclint/_0015_ ), .Z(\myclint/_0473_ ) );
BUF_X1 \myclint/_1040_ ( .A(\myclint/_0016_ ), .Z(\myclint/_0474_ ) );
BUF_X1 \myclint/_1041_ ( .A(\myclint/_0017_ ), .Z(\myclint/_0475_ ) );
BUF_X1 \myclint/_1042_ ( .A(\myclint/_0018_ ), .Z(\myclint/_0476_ ) );
BUF_X1 \myclint/_1043_ ( .A(\myclint/_0019_ ), .Z(\myclint/_0477_ ) );
BUF_X1 \myclint/_1044_ ( .A(\myclint/_0020_ ), .Z(\myclint/_0478_ ) );
BUF_X1 \myclint/_1045_ ( .A(\myclint/_0021_ ), .Z(\myclint/_0479_ ) );
BUF_X1 \myclint/_1046_ ( .A(\myclint/_0022_ ), .Z(\myclint/_0480_ ) );
BUF_X1 \myclint/_1047_ ( .A(\myclint/_0023_ ), .Z(\myclint/_0481_ ) );
BUF_X1 \myclint/_1048_ ( .A(\myclint/_0024_ ), .Z(\myclint/_0482_ ) );
BUF_X1 \myclint/_1049_ ( .A(\myclint/_0025_ ), .Z(\myclint/_0483_ ) );
BUF_X1 \myclint/_1050_ ( .A(\myclint/_0026_ ), .Z(\myclint/_0484_ ) );
BUF_X1 \myclint/_1051_ ( .A(\myclint/_0027_ ), .Z(\myclint/_0485_ ) );
BUF_X1 \myclint/_1052_ ( .A(\myclint/_0028_ ), .Z(\myclint/_0486_ ) );
BUF_X1 \myclint/_1053_ ( .A(\myclint/_0029_ ), .Z(\myclint/_0487_ ) );
BUF_X1 \myclint/_1054_ ( .A(\myclint/_0030_ ), .Z(\myclint/_0488_ ) );
BUF_X1 \myclint/_1055_ ( .A(\myclint/_0031_ ), .Z(\myclint/_0489_ ) );
BUF_X1 \myclint/_1056_ ( .A(\myclint/_0032_ ), .Z(\myclint/_0490_ ) );
BUF_X1 \myclint/_1057_ ( .A(\myclint/_0033_ ), .Z(\myclint/_0491_ ) );
BUF_X1 \myclint/_1058_ ( .A(\myclint/_0034_ ), .Z(\myclint/_0492_ ) );
BUF_X1 \myclint/_1059_ ( .A(\myclint/_0035_ ), .Z(\myclint/_0493_ ) );
BUF_X1 \myclint/_1060_ ( .A(\myclint/_0036_ ), .Z(\myclint/_0494_ ) );
BUF_X1 \myclint/_1061_ ( .A(\myclint/_0037_ ), .Z(\myclint/_0495_ ) );
BUF_X1 \myclint/_1062_ ( .A(\myclint/_0038_ ), .Z(\myclint/_0496_ ) );
BUF_X1 \myclint/_1063_ ( .A(\myclint/_0039_ ), .Z(\myclint/_0497_ ) );
BUF_X1 \myclint/_1064_ ( .A(\myclint/_0040_ ), .Z(\myclint/_0498_ ) );
BUF_X1 \myclint/_1065_ ( .A(\myclint/_0041_ ), .Z(\myclint/_0499_ ) );
BUF_X1 \myclint/_1066_ ( .A(\myclint/_0042_ ), .Z(\myclint/_0500_ ) );
BUF_X1 \myclint/_1067_ ( .A(\myclint/_0043_ ), .Z(\myclint/_0501_ ) );
BUF_X1 \myclint/_1068_ ( .A(\myclint/_0044_ ), .Z(\myclint/_0502_ ) );
BUF_X1 \myclint/_1069_ ( .A(\myclint/_0045_ ), .Z(\myclint/_0503_ ) );
BUF_X1 \myclint/_1070_ ( .A(\myclint/_0046_ ), .Z(\myclint/_0504_ ) );
BUF_X1 \myclint/_1071_ ( .A(\myclint/_0047_ ), .Z(\myclint/_0505_ ) );
BUF_X1 \myclint/_1072_ ( .A(\myclint/_0048_ ), .Z(\myclint/_0506_ ) );
BUF_X1 \myclint/_1073_ ( .A(\myclint/_0049_ ), .Z(\myclint/_0507_ ) );
BUF_X1 \myclint/_1074_ ( .A(\myclint/_0050_ ), .Z(\myclint/_0508_ ) );
BUF_X1 \myclint/_1075_ ( .A(\myclint/_0051_ ), .Z(\myclint/_0509_ ) );
BUF_X1 \myclint/_1076_ ( .A(\myclint/_0052_ ), .Z(\myclint/_0510_ ) );
BUF_X1 \myclint/_1077_ ( .A(\myclint/_0053_ ), .Z(\myclint/_0511_ ) );
BUF_X1 \myclint/_1078_ ( .A(\myclint/_0054_ ), .Z(\myclint/_0512_ ) );
BUF_X1 \myclint/_1079_ ( .A(\myclint/_0055_ ), .Z(\myclint/_0513_ ) );
BUF_X1 \myclint/_1080_ ( .A(\myclint/_0056_ ), .Z(\myclint/_0514_ ) );
BUF_X1 \myclint/_1081_ ( .A(\myclint/_0057_ ), .Z(\myclint/_0515_ ) );
BUF_X1 \myclint/_1082_ ( .A(\myclint/_0058_ ), .Z(\myclint/_0516_ ) );
BUF_X1 \myclint/_1083_ ( .A(\myclint/_0059_ ), .Z(\myclint/_0517_ ) );
BUF_X1 \myclint/_1084_ ( .A(\myclint/_0060_ ), .Z(\myclint/_0518_ ) );
BUF_X1 \myclint/_1085_ ( .A(\myclint/_0061_ ), .Z(\myclint/_0519_ ) );
BUF_X1 \myclint/_1086_ ( .A(\myclint/_0062_ ), .Z(\myclint/_0520_ ) );
BUF_X1 \myclint/_1087_ ( .A(\myclint/_0063_ ), .Z(\myclint/_0521_ ) );
BUF_X1 \myclint/_1088_ ( .A(\myclint/_0064_ ), .Z(\myclint/_0522_ ) );
BUF_X1 \myclint/_1089_ ( .A(\myclint/_0065_ ), .Z(\myclint/_0523_ ) );
BUF_X1 \myclint/_1090_ ( .A(\myclint/_0066_ ), .Z(\myclint/_0524_ ) );
BUF_X1 \myclint/_1091_ ( .A(\myclint/_0067_ ), .Z(\myclint/_0525_ ) );
AND2_X1 \mycsreg/_0932_ ( .A1(\mycsreg/_0590_ ), .A2(\mycsreg/_0589_ ), .ZN(\mycsreg/_0256_ ) );
INV_X1 \mycsreg/_0933_ ( .A(\mycsreg/_0256_ ), .ZN(\mycsreg/_0257_ ) );
NOR3_X1 \mycsreg/_0934_ ( .A1(\mycsreg/_0257_ ), .A2(\mycsreg/_0581_ ), .A3(\mycsreg/_0580_ ), .ZN(\mycsreg/_0258_ ) );
CLKBUF_X2 \mycsreg/_0935_ ( .A(\mycsreg/_0258_ ), .Z(\mycsreg/_0259_ ) );
INV_X16 \mycsreg/_0936_ ( .A(\mycsreg/_0585_ ), .ZN(\mycsreg/_0260_ ) );
NAND2_X1 \mycsreg/_0937_ ( .A1(\mycsreg/_0260_ ), .A2(\mycsreg/_0587_ ), .ZN(\mycsreg/_0261_ ) );
NOR3_X4 \mycsreg/_0938_ ( .A1(\mycsreg/_0261_ ), .A2(\mycsreg/_0588_ ), .A3(\mycsreg/_0586_ ), .ZN(\mycsreg/_0262_ ) );
BUF_X2 \mycsreg/_0939_ ( .A(\mycsreg/_0262_ ), .Z(\mycsreg/_0263_ ) );
NOR2_X1 \mycsreg/_0940_ ( .A1(\mycsreg/_0584_ ), .A2(\mycsreg/_0583_ ), .ZN(\mycsreg/_0264_ ) );
INV_X1 \mycsreg/_0941_ ( .A(\mycsreg/_0264_ ), .ZN(\mycsreg/_0265_ ) );
INV_X1 \mycsreg/_0942_ ( .A(\mycsreg/_0579_ ), .ZN(\mycsreg/_0266_ ) );
NOR3_X2 \mycsreg/_0943_ ( .A1(\mycsreg/_0265_ ), .A2(\mycsreg/_0582_ ), .A3(\mycsreg/_0266_ ), .ZN(\mycsreg/_0267_ ) );
AND4_X1 \mycsreg/_0944_ ( .A1(\mycsreg/_0064_ ), .A2(\mycsreg/_0259_ ), .A3(\mycsreg/_0263_ ), .A4(\mycsreg/_0267_ ), .ZN(\mycsreg/_0268_ ) );
AND3_X1 \mycsreg/_0945_ ( .A1(\mycsreg/_0264_ ), .A2(\mycsreg/_0582_ ), .A3(\mycsreg/_0266_ ), .ZN(\mycsreg/_0269_ ) );
BUF_X4 \mycsreg/_0946_ ( .A(\mycsreg/_0269_ ), .Z(\mycsreg/_0270_ ) );
BUF_X4 \mycsreg/_0947_ ( .A(\mycsreg/_0270_ ), .Z(\mycsreg/_0271_ ) );
BUF_X4 \mycsreg/_0948_ ( .A(\mycsreg/_0271_ ), .Z(\mycsreg/_0272_ ) );
AND4_X1 \mycsreg/_0949_ ( .A1(\mycsreg/_0581_ ), .A2(\mycsreg/_0256_ ), .A3(\mycsreg/_0580_ ), .A4(\mycsreg/_0585_ ), .ZN(\mycsreg/_0273_ ) );
NOR3_X1 \mycsreg/_0950_ ( .A1(\mycsreg/_0588_ ), .A2(\mycsreg/_0587_ ), .A3(\mycsreg/_0586_ ), .ZN(\mycsreg/_0274_ ) );
AND2_X2 \mycsreg/_0951_ ( .A1(\mycsreg/_0273_ ), .A2(\mycsreg/_0274_ ), .ZN(\mycsreg/_0275_ ) );
AOI21_X1 \mycsreg/_0952_ ( .A(\mycsreg/_0268_ ), .B1(\mycsreg/_0272_ ), .B2(\mycsreg/_0275_ ), .ZN(\mycsreg/_0276_ ) );
BUF_X8 \mycsreg/_0953_ ( .A(\mycsreg/_0258_ ), .Z(\mycsreg/_0277_ ) );
BUF_X4 \mycsreg/_0954_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0278_ ) );
AND2_X1 \mycsreg/_0955_ ( .A1(\mycsreg/_0274_ ), .A2(\mycsreg/_0260_ ), .ZN(\mycsreg/_0279_ ) );
BUF_X4 \mycsreg/_0956_ ( .A(\mycsreg/_0279_ ), .Z(\mycsreg/_0280_ ) );
BUF_X4 \mycsreg/_0957_ ( .A(\mycsreg/_0280_ ), .Z(\mycsreg/_0281_ ) );
INV_X1 \mycsreg/_0958_ ( .A(\mycsreg/_0583_ ), .ZN(\mycsreg/_0282_ ) );
NOR4_X2 \mycsreg/_0959_ ( .A1(\mycsreg/_0282_ ), .A2(\mycsreg/_0266_ ), .A3(\mycsreg/_0584_ ), .A4(\mycsreg/_0582_ ), .ZN(\mycsreg/_0283_ ) );
BUF_X4 \mycsreg/_0960_ ( .A(\mycsreg/_0283_ ), .Z(\mycsreg/_0284_ ) );
NAND4_X1 \mycsreg/_0961_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0032_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0285_ ) );
BUF_X4 \mycsreg/_0962_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0286_ ) );
BUF_X4 \mycsreg/_0963_ ( .A(\mycsreg/_0280_ ), .Z(\mycsreg/_0287_ ) );
NOR4_X2 \mycsreg/_0964_ ( .A1(\mycsreg/_0584_ ), .A2(\mycsreg/_0583_ ), .A3(\mycsreg/_0582_ ), .A4(\mycsreg/_0579_ ), .ZN(\mycsreg/_0288_ ) );
BUF_X4 \mycsreg/_0965_ ( .A(\mycsreg/_0288_ ), .Z(\mycsreg/_0289_ ) );
NAND4_X1 \mycsreg/_0966_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0000_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0290_ ) );
BUF_X4 \mycsreg/_0967_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0291_ ) );
BUF_X4 \mycsreg/_0968_ ( .A(\mycsreg/_0262_ ), .Z(\mycsreg/_0292_ ) );
NAND4_X1 \mycsreg/_0969_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0096_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0293_ ) );
AND3_X1 \mycsreg/_0970_ ( .A1(\mycsreg/_0285_ ), .A2(\mycsreg/_0290_ ), .A3(\mycsreg/_0293_ ), .ZN(\mycsreg/_0294_ ) );
NAND2_X1 \mycsreg/_0971_ ( .A1(\mycsreg/_0276_ ), .A2(\mycsreg/_0294_ ), .ZN(\mycsreg/_0591_ ) );
BUF_X4 \mycsreg/_0972_ ( .A(\mycsreg/_0278_ ), .Z(\mycsreg/_0295_ ) );
BUF_X4 \mycsreg/_0973_ ( .A(\mycsreg/_0267_ ), .Z(\mycsreg/_0296_ ) );
BUF_X4 \mycsreg/_0974_ ( .A(\mycsreg/_0296_ ), .Z(\mycsreg/_0297_ ) );
BUF_X4 \mycsreg/_0975_ ( .A(\mycsreg/_0262_ ), .Z(\mycsreg/_0298_ ) );
BUF_X4 \mycsreg/_0976_ ( .A(\mycsreg/_0298_ ), .Z(\mycsreg/_0299_ ) );
NAND4_X1 \mycsreg/_0977_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0297_ ), .A3(\mycsreg/_0075_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0300_ ) );
BUF_X4 \mycsreg/_0978_ ( .A(\mycsreg/_0286_ ), .Z(\mycsreg/_0301_ ) );
BUF_X4 \mycsreg/_0979_ ( .A(\mycsreg/_0287_ ), .Z(\mycsreg/_0302_ ) );
NAND4_X1 \mycsreg/_0980_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0043_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0303_ ) );
BUF_X4 \mycsreg/_0981_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0304_ ) );
BUF_X4 \mycsreg/_0982_ ( .A(\mycsreg/_0304_ ), .Z(\mycsreg/_0305_ ) );
NAND4_X1 \mycsreg/_0983_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0107_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0306_ ) );
NAND4_X1 \mycsreg/_0984_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0011_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0307_ ) );
NAND4_X1 \mycsreg/_0985_ ( .A1(\mycsreg/_0300_ ), .A2(\mycsreg/_0303_ ), .A3(\mycsreg/_0306_ ), .A4(\mycsreg/_0307_ ), .ZN(\mycsreg/_0602_ ) );
BUF_X4 \mycsreg/_0986_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0308_ ) );
BUF_X4 \mycsreg/_0987_ ( .A(\mycsreg/_0270_ ), .Z(\mycsreg/_0309_ ) );
BUF_X4 \mycsreg/_0988_ ( .A(\mycsreg/_0262_ ), .Z(\mycsreg/_0310_ ) );
NAND4_X1 \mycsreg/_0989_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0118_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0311_ ) );
BUF_X4 \mycsreg/_0990_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0312_ ) );
BUF_X4 \mycsreg/_0991_ ( .A(\mycsreg/_0267_ ), .Z(\mycsreg/_0313_ ) );
NAND4_X1 \mycsreg/_0992_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0086_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0314_ ) );
BUF_X4 \mycsreg/_0993_ ( .A(\mycsreg/_0280_ ), .Z(\mycsreg/_0315_ ) );
BUF_X4 \mycsreg/_0994_ ( .A(\mycsreg/_0283_ ), .Z(\mycsreg/_0316_ ) );
NAND4_X1 \mycsreg/_0995_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0054_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0317_ ) );
AND3_X1 \mycsreg/_0996_ ( .A1(\mycsreg/_0311_ ), .A2(\mycsreg/_0314_ ), .A3(\mycsreg/_0317_ ), .ZN(\mycsreg/_0318_ ) );
AND2_X1 \mycsreg/_0997_ ( .A1(\mycsreg/_0275_ ), .A2(\mycsreg/_0270_ ), .ZN(\mycsreg/_0319_ ) );
INV_X1 \mycsreg/_0998_ ( .A(\mycsreg/_0319_ ), .ZN(\mycsreg/_0320_ ) );
BUF_X4 \mycsreg/_0999_ ( .A(\mycsreg/_0320_ ), .Z(\mycsreg/_0321_ ) );
BUF_X4 \mycsreg/_1000_ ( .A(\mycsreg/_0289_ ), .Z(\mycsreg/_0322_ ) );
NAND4_X1 \mycsreg/_1001_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0022_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0323_ ) );
NAND3_X1 \mycsreg/_1002_ ( .A1(\mycsreg/_0318_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0323_ ), .ZN(\mycsreg/_0613_ ) );
NAND4_X1 \mycsreg/_1003_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0057_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0324_ ) );
NAND4_X1 \mycsreg/_1004_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0025_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0325_ ) );
NAND4_X1 \mycsreg/_1005_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0121_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0326_ ) );
AND3_X1 \mycsreg/_1006_ ( .A1(\mycsreg/_0324_ ), .A2(\mycsreg/_0325_ ), .A3(\mycsreg/_0326_ ), .ZN(\mycsreg/_0327_ ) );
AND2_X1 \mycsreg/_1007_ ( .A1(\mycsreg/_0275_ ), .A2(\mycsreg/_0267_ ), .ZN(\mycsreg/_0328_ ) );
INV_X1 \mycsreg/_1008_ ( .A(\mycsreg/_0328_ ), .ZN(\mycsreg/_0329_ ) );
BUF_X4 \mycsreg/_1009_ ( .A(\mycsreg/_0329_ ), .Z(\mycsreg/_0330_ ) );
NAND4_X1 \mycsreg/_1010_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0297_ ), .A3(\mycsreg/_0089_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0331_ ) );
NAND3_X1 \mycsreg/_1011_ ( .A1(\mycsreg/_0327_ ), .A2(\mycsreg/_0330_ ), .A3(\mycsreg/_0331_ ), .ZN(\mycsreg/_0616_ ) );
AND4_X1 \mycsreg/_1012_ ( .A1(\mycsreg/_0122_ ), .A2(\mycsreg/_0259_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0332_ ) );
AOI21_X1 \mycsreg/_1013_ ( .A(\mycsreg/_0332_ ), .B1(\mycsreg/_0275_ ), .B2(\mycsreg/_0297_ ), .ZN(\mycsreg/_0333_ ) );
NAND4_X1 \mycsreg/_1014_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0090_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0334_ ) );
NAND4_X1 \mycsreg/_1015_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0058_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0335_ ) );
NAND4_X1 \mycsreg/_1016_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0026_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0336_ ) );
AND3_X1 \mycsreg/_1017_ ( .A1(\mycsreg/_0334_ ), .A2(\mycsreg/_0335_ ), .A3(\mycsreg/_0336_ ), .ZN(\mycsreg/_0337_ ) );
NAND2_X1 \mycsreg/_1018_ ( .A1(\mycsreg/_0333_ ), .A2(\mycsreg/_0337_ ), .ZN(\mycsreg/_0617_ ) );
BUF_X4 \mycsreg/_1019_ ( .A(\mycsreg/_0262_ ), .Z(\mycsreg/_0338_ ) );
NAND4_X1 \mycsreg/_1020_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0123_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0339_ ) );
NAND4_X1 \mycsreg/_1021_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0091_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0340_ ) );
NAND4_X1 \mycsreg/_1022_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0059_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0341_ ) );
AND3_X1 \mycsreg/_1023_ ( .A1(\mycsreg/_0339_ ), .A2(\mycsreg/_0340_ ), .A3(\mycsreg/_0341_ ), .ZN(\mycsreg/_0342_ ) );
NAND4_X1 \mycsreg/_1024_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0027_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0343_ ) );
NAND3_X1 \mycsreg/_1025_ ( .A1(\mycsreg/_0342_ ), .A2(\mycsreg/_0330_ ), .A3(\mycsreg/_0343_ ), .ZN(\mycsreg/_0618_ ) );
BUF_X2 \mycsreg/_1026_ ( .A(\mycsreg/_0280_ ), .Z(\mycsreg/_0344_ ) );
BUF_X2 \mycsreg/_1027_ ( .A(\mycsreg/_0288_ ), .Z(\mycsreg/_0345_ ) );
AND4_X2 \mycsreg/_1028_ ( .A1(\mycsreg/_0028_ ), .A2(\mycsreg/_0259_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0346_ ) );
AOI21_X1 \mycsreg/_1029_ ( .A(\mycsreg/_0346_ ), .B1(\mycsreg/_0275_ ), .B2(\mycsreg/_0297_ ), .ZN(\mycsreg/_0347_ ) );
NAND4_X1 \mycsreg/_1030_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0124_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0348_ ) );
NAND4_X1 \mycsreg/_1031_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0092_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0349_ ) );
NAND4_X1 \mycsreg/_1032_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0060_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0350_ ) );
AND3_X1 \mycsreg/_1033_ ( .A1(\mycsreg/_0348_ ), .A2(\mycsreg/_0349_ ), .A3(\mycsreg/_0350_ ), .ZN(\mycsreg/_0351_ ) );
NAND2_X1 \mycsreg/_1034_ ( .A1(\mycsreg/_0347_ ), .A2(\mycsreg/_0351_ ), .ZN(\mycsreg/_0619_ ) );
NAND4_X1 \mycsreg/_1035_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0297_ ), .A3(\mycsreg/_0093_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0352_ ) );
NAND4_X1 \mycsreg/_1036_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0029_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0353_ ) );
NAND4_X1 \mycsreg/_1037_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0125_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0354_ ) );
NAND4_X1 \mycsreg/_1038_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0061_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0355_ ) );
NAND4_X1 \mycsreg/_1039_ ( .A1(\mycsreg/_0352_ ), .A2(\mycsreg/_0353_ ), .A3(\mycsreg/_0354_ ), .A4(\mycsreg/_0355_ ), .ZN(\mycsreg/_0620_ ) );
NAND4_X1 \mycsreg/_1040_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0094_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0356_ ) );
BUF_X4 \mycsreg/_1041_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0357_ ) );
BUF_X4 \mycsreg/_1042_ ( .A(\mycsreg/_0280_ ), .Z(\mycsreg/_0358_ ) );
BUF_X2 \mycsreg/_1043_ ( .A(\mycsreg/_0283_ ), .Z(\mycsreg/_0359_ ) );
NAND4_X1 \mycsreg/_1044_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0062_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0360_ ) );
BUF_X4 \mycsreg/_1045_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0361_ ) );
NAND4_X1 \mycsreg/_1046_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0126_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0362_ ) );
BUF_X4 \mycsreg/_1047_ ( .A(\mycsreg/_0277_ ), .Z(\mycsreg/_0363_ ) );
NAND4_X1 \mycsreg/_1048_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0030_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0364_ ) );
AND4_X1 \mycsreg/_1049_ ( .A1(\mycsreg/_0356_ ), .A2(\mycsreg/_0360_ ), .A3(\mycsreg/_0362_ ), .A4(\mycsreg/_0364_ ), .ZN(\mycsreg/_0365_ ) );
NAND3_X1 \mycsreg/_1050_ ( .A1(\mycsreg/_0365_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0330_ ), .ZN(\mycsreg/_0621_ ) );
NAND4_X1 \mycsreg/_1051_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0127_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0366_ ) );
NAND4_X1 \mycsreg/_1052_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0095_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0367_ ) );
NAND4_X1 \mycsreg/_1053_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0063_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0368_ ) );
AND3_X1 \mycsreg/_1054_ ( .A1(\mycsreg/_0366_ ), .A2(\mycsreg/_0367_ ), .A3(\mycsreg/_0368_ ), .ZN(\mycsreg/_0369_ ) );
NAND4_X1 \mycsreg/_1055_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0031_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0370_ ) );
NAND3_X1 \mycsreg/_1056_ ( .A1(\mycsreg/_0369_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0370_ ), .ZN(\mycsreg/_0622_ ) );
AND4_X2 \mycsreg/_1057_ ( .A1(\mycsreg/_0001_ ), .A2(\mycsreg/_0259_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0371_ ) );
AOI21_X1 \mycsreg/_1058_ ( .A(\mycsreg/_0371_ ), .B1(\mycsreg/_0272_ ), .B2(\mycsreg/_0275_ ), .ZN(\mycsreg/_0372_ ) );
NAND4_X1 \mycsreg/_1059_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0097_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0373_ ) );
NAND4_X1 \mycsreg/_1060_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0065_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0374_ ) );
NAND4_X1 \mycsreg/_1061_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0033_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0375_ ) );
AND3_X1 \mycsreg/_1062_ ( .A1(\mycsreg/_0373_ ), .A2(\mycsreg/_0374_ ), .A3(\mycsreg/_0375_ ), .ZN(\mycsreg/_0376_ ) );
NAND2_X1 \mycsreg/_1063_ ( .A1(\mycsreg/_0372_ ), .A2(\mycsreg/_0376_ ), .ZN(\mycsreg/_0592_ ) );
NAND4_X1 \mycsreg/_1064_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0066_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0377_ ) );
NAND4_X1 \mycsreg/_1065_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0034_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0378_ ) );
NAND4_X1 \mycsreg/_1066_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0098_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0379_ ) );
NAND4_X1 \mycsreg/_1067_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0002_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0380_ ) );
AND4_X1 \mycsreg/_1068_ ( .A1(\mycsreg/_0377_ ), .A2(\mycsreg/_0378_ ), .A3(\mycsreg/_0379_ ), .A4(\mycsreg/_0380_ ), .ZN(\mycsreg/_0381_ ) );
NAND3_X1 \mycsreg/_1069_ ( .A1(\mycsreg/_0381_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0330_ ), .ZN(\mycsreg/_0593_ ) );
NAND4_X1 \mycsreg/_1070_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0067_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0382_ ) );
NAND4_X1 \mycsreg/_1071_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0035_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0383_ ) );
NAND4_X1 \mycsreg/_1072_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0099_ ), .A3(\mycsreg/_0270_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0384_ ) );
NAND4_X1 \mycsreg/_1073_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0003_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0385_ ) );
AND4_X1 \mycsreg/_1074_ ( .A1(\mycsreg/_0382_ ), .A2(\mycsreg/_0383_ ), .A3(\mycsreg/_0384_ ), .A4(\mycsreg/_0385_ ), .ZN(\mycsreg/_0386_ ) );
NAND3_X1 \mycsreg/_1075_ ( .A1(\mycsreg/_0386_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0330_ ), .ZN(\mycsreg/_0594_ ) );
NAND4_X1 \mycsreg/_1076_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0036_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0387_ ) );
NAND4_X1 \mycsreg/_1077_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0004_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0388_ ) );
NAND4_X1 \mycsreg/_1078_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0100_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0389_ ) );
AND3_X1 \mycsreg/_1079_ ( .A1(\mycsreg/_0387_ ), .A2(\mycsreg/_0388_ ), .A3(\mycsreg/_0389_ ), .ZN(\mycsreg/_0390_ ) );
NAND4_X1 \mycsreg/_1080_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0297_ ), .A3(\mycsreg/_0068_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0391_ ) );
NAND3_X1 \mycsreg/_1081_ ( .A1(\mycsreg/_0390_ ), .A2(\mycsreg/_0330_ ), .A3(\mycsreg/_0391_ ), .ZN(\mycsreg/_0595_ ) );
NAND4_X1 \mycsreg/_1082_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0101_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0392_ ) );
NAND4_X1 \mycsreg/_1083_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0005_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0393_ ) );
NAND4_X1 \mycsreg/_1084_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0267_ ), .A3(\mycsreg/_0069_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0394_ ) );
NAND4_X1 \mycsreg/_1085_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0037_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0283_ ), .ZN(\mycsreg/_0395_ ) );
AND4_X1 \mycsreg/_1086_ ( .A1(\mycsreg/_0392_ ), .A2(\mycsreg/_0393_ ), .A3(\mycsreg/_0394_ ), .A4(\mycsreg/_0395_ ), .ZN(\mycsreg/_0396_ ) );
NAND3_X1 \mycsreg/_1087_ ( .A1(\mycsreg/_0396_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0330_ ), .ZN(\mycsreg/_0596_ ) );
NAND4_X1 \mycsreg/_1088_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0006_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0397_ ) );
NAND4_X1 \mycsreg/_1089_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0102_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0398_ ) );
NAND4_X1 \mycsreg/_1090_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0070_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0399_ ) );
AND3_X1 \mycsreg/_1091_ ( .A1(\mycsreg/_0397_ ), .A2(\mycsreg/_0398_ ), .A3(\mycsreg/_0399_ ), .ZN(\mycsreg/_0400_ ) );
NAND4_X1 \mycsreg/_1092_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0038_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0401_ ) );
NAND3_X1 \mycsreg/_1093_ ( .A1(\mycsreg/_0400_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0401_ ), .ZN(\mycsreg/_0597_ ) );
NAND4_X1 \mycsreg/_1094_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0267_ ), .A3(\mycsreg/_0071_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0402_ ) );
NAND4_X1 \mycsreg/_1095_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0039_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0403_ ) );
NAND4_X1 \mycsreg/_1096_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0103_ ), .A3(\mycsreg/_0270_ ), .A4(\mycsreg/_0262_ ), .ZN(\mycsreg/_0404_ ) );
NAND4_X1 \mycsreg/_1097_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0007_ ), .A3(\mycsreg/_0280_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0405_ ) );
AND4_X1 \mycsreg/_1098_ ( .A1(\mycsreg/_0402_ ), .A2(\mycsreg/_0403_ ), .A3(\mycsreg/_0404_ ), .A4(\mycsreg/_0405_ ), .ZN(\mycsreg/_0406_ ) );
NAND3_X1 \mycsreg/_1099_ ( .A1(\mycsreg/_0406_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0329_ ), .ZN(\mycsreg/_0598_ ) );
NAND4_X1 \mycsreg/_1100_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0267_ ), .A3(\mycsreg/_0072_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0407_ ) );
NAND4_X1 \mycsreg/_1101_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0040_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0408_ ) );
NAND4_X1 \mycsreg/_1102_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0104_ ), .A3(\mycsreg/_0270_ ), .A4(\mycsreg/_0262_ ), .ZN(\mycsreg/_0409_ ) );
NAND4_X1 \mycsreg/_1103_ ( .A1(\mycsreg/_0259_ ), .A2(\mycsreg/_0008_ ), .A3(\mycsreg/_0280_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0410_ ) );
AND4_X1 \mycsreg/_1104_ ( .A1(\mycsreg/_0407_ ), .A2(\mycsreg/_0408_ ), .A3(\mycsreg/_0409_ ), .A4(\mycsreg/_0410_ ), .ZN(\mycsreg/_0411_ ) );
NAND3_X1 \mycsreg/_1105_ ( .A1(\mycsreg/_0411_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0329_ ), .ZN(\mycsreg/_0599_ ) );
NAND4_X1 \mycsreg/_1106_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0105_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0412_ ) );
NAND4_X1 \mycsreg/_1107_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0073_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0413_ ) );
NAND4_X1 \mycsreg/_1108_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0041_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0414_ ) );
AND3_X1 \mycsreg/_1109_ ( .A1(\mycsreg/_0412_ ), .A2(\mycsreg/_0413_ ), .A3(\mycsreg/_0414_ ), .ZN(\mycsreg/_0415_ ) );
NAND4_X1 \mycsreg/_1110_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0009_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0416_ ) );
NAND3_X1 \mycsreg/_1111_ ( .A1(\mycsreg/_0415_ ), .A2(\mycsreg/_0321_ ), .A3(\mycsreg/_0416_ ), .ZN(\mycsreg/_0600_ ) );
AND4_X2 \mycsreg/_1112_ ( .A1(\mycsreg/_0010_ ), .A2(\mycsreg/_0259_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0417_ ) );
AOI21_X1 \mycsreg/_1113_ ( .A(\mycsreg/_0417_ ), .B1(\mycsreg/_0272_ ), .B2(\mycsreg/_0275_ ), .ZN(\mycsreg/_0418_ ) );
NAND4_X1 \mycsreg/_1114_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0106_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0419_ ) );
NAND4_X1 \mycsreg/_1115_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0074_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0420_ ) );
NAND4_X1 \mycsreg/_1116_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0042_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0421_ ) );
AND3_X1 \mycsreg/_1117_ ( .A1(\mycsreg/_0419_ ), .A2(\mycsreg/_0420_ ), .A3(\mycsreg/_0421_ ), .ZN(\mycsreg/_0422_ ) );
NAND2_X1 \mycsreg/_1118_ ( .A1(\mycsreg/_0418_ ), .A2(\mycsreg/_0422_ ), .ZN(\mycsreg/_0601_ ) );
NAND4_X1 \mycsreg/_1119_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0267_ ), .A3(\mycsreg/_0076_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0423_ ) );
NAND4_X1 \mycsreg/_1120_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0044_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0424_ ) );
NAND4_X1 \mycsreg/_1121_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0108_ ), .A3(\mycsreg/_0270_ ), .A4(\mycsreg/_0262_ ), .ZN(\mycsreg/_0425_ ) );
NAND4_X1 \mycsreg/_1122_ ( .A1(\mycsreg/_0259_ ), .A2(\mycsreg/_0012_ ), .A3(\mycsreg/_0280_ ), .A4(\mycsreg/_0288_ ), .ZN(\mycsreg/_0426_ ) );
AND4_X2 \mycsreg/_1123_ ( .A1(\mycsreg/_0423_ ), .A2(\mycsreg/_0424_ ), .A3(\mycsreg/_0425_ ), .A4(\mycsreg/_0426_ ), .ZN(\mycsreg/_0427_ ) );
NAND3_X1 \mycsreg/_1124_ ( .A1(\mycsreg/_0427_ ), .A2(\mycsreg/_0320_ ), .A3(\mycsreg/_0329_ ), .ZN(\mycsreg/_0603_ ) );
AND4_X1 \mycsreg/_1125_ ( .A1(\mycsreg/_0045_ ), .A2(\mycsreg/_0259_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0428_ ) );
AOI21_X1 \mycsreg/_1126_ ( .A(\mycsreg/_0428_ ), .B1(\mycsreg/_0275_ ), .B2(\mycsreg/_0297_ ), .ZN(\mycsreg/_0429_ ) );
NAND4_X1 \mycsreg/_1127_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0013_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0430_ ) );
NAND4_X1 \mycsreg/_1128_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0109_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0431_ ) );
NAND4_X1 \mycsreg/_1129_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0077_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0432_ ) );
AND3_X1 \mycsreg/_1130_ ( .A1(\mycsreg/_0430_ ), .A2(\mycsreg/_0431_ ), .A3(\mycsreg/_0432_ ), .ZN(\mycsreg/_0433_ ) );
NAND2_X1 \mycsreg/_1131_ ( .A1(\mycsreg/_0429_ ), .A2(\mycsreg/_0433_ ), .ZN(\mycsreg/_0604_ ) );
NAND4_X1 \mycsreg/_1132_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0267_ ), .A3(\mycsreg/_0078_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0434_ ) );
NAND4_X1 \mycsreg/_1133_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0046_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0435_ ) );
NAND4_X1 \mycsreg/_1134_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0110_ ), .A3(\mycsreg/_0270_ ), .A4(\mycsreg/_0262_ ), .ZN(\mycsreg/_0436_ ) );
NAND4_X1 \mycsreg/_1135_ ( .A1(\mycsreg/_0259_ ), .A2(\mycsreg/_0014_ ), .A3(\mycsreg/_0280_ ), .A4(\mycsreg/_0288_ ), .ZN(\mycsreg/_0437_ ) );
AND4_X1 \mycsreg/_1136_ ( .A1(\mycsreg/_0434_ ), .A2(\mycsreg/_0435_ ), .A3(\mycsreg/_0436_ ), .A4(\mycsreg/_0437_ ), .ZN(\mycsreg/_0438_ ) );
NAND3_X1 \mycsreg/_1137_ ( .A1(\mycsreg/_0438_ ), .A2(\mycsreg/_0320_ ), .A3(\mycsreg/_0329_ ), .ZN(\mycsreg/_0605_ ) );
NAND4_X1 \mycsreg/_1138_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0111_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0439_ ) );
NAND4_X1 \mycsreg/_1139_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0015_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0440_ ) );
NAND4_X1 \mycsreg/_1140_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0297_ ), .A3(\mycsreg/_0079_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0441_ ) );
NAND4_X1 \mycsreg/_1141_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0047_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0442_ ) );
NAND4_X1 \mycsreg/_1142_ ( .A1(\mycsreg/_0439_ ), .A2(\mycsreg/_0440_ ), .A3(\mycsreg/_0441_ ), .A4(\mycsreg/_0442_ ), .ZN(\mycsreg/_0606_ ) );
NAND4_X1 \mycsreg/_1143_ ( .A1(\mycsreg/_0357_ ), .A2(\mycsreg/_0267_ ), .A3(\mycsreg/_0080_ ), .A4(\mycsreg/_0263_ ), .ZN(\mycsreg/_0443_ ) );
NAND4_X1 \mycsreg/_1144_ ( .A1(\mycsreg/_0361_ ), .A2(\mycsreg/_0048_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0444_ ) );
NAND4_X1 \mycsreg/_1145_ ( .A1(\mycsreg/_0363_ ), .A2(\mycsreg/_0112_ ), .A3(\mycsreg/_0270_ ), .A4(\mycsreg/_0262_ ), .ZN(\mycsreg/_0445_ ) );
NAND4_X1 \mycsreg/_1146_ ( .A1(\mycsreg/_0259_ ), .A2(\mycsreg/_0016_ ), .A3(\mycsreg/_0280_ ), .A4(\mycsreg/_0288_ ), .ZN(\mycsreg/_0446_ ) );
AND4_X1 \mycsreg/_1147_ ( .A1(\mycsreg/_0443_ ), .A2(\mycsreg/_0444_ ), .A3(\mycsreg/_0445_ ), .A4(\mycsreg/_0446_ ), .ZN(\mycsreg/_0447_ ) );
NAND3_X1 \mycsreg/_1148_ ( .A1(\mycsreg/_0447_ ), .A2(\mycsreg/_0320_ ), .A3(\mycsreg/_0329_ ), .ZN(\mycsreg/_0607_ ) );
NAND4_X1 \mycsreg/_1149_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0113_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0448_ ) );
NAND4_X1 \mycsreg/_1150_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0017_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0449_ ) );
NAND4_X1 \mycsreg/_1151_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0081_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0450_ ) );
NAND4_X1 \mycsreg/_1152_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0049_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0451_ ) );
NAND4_X1 \mycsreg/_1153_ ( .A1(\mycsreg/_0448_ ), .A2(\mycsreg/_0449_ ), .A3(\mycsreg/_0450_ ), .A4(\mycsreg/_0451_ ), .ZN(\mycsreg/_0608_ ) );
NAND4_X1 \mycsreg/_1154_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0297_ ), .A3(\mycsreg/_0082_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0452_ ) );
NAND4_X1 \mycsreg/_1155_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0018_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0453_ ) );
NAND4_X1 \mycsreg/_1156_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0114_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0454_ ) );
NAND4_X1 \mycsreg/_1157_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0050_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0455_ ) );
NAND4_X1 \mycsreg/_1158_ ( .A1(\mycsreg/_0452_ ), .A2(\mycsreg/_0453_ ), .A3(\mycsreg/_0454_ ), .A4(\mycsreg/_0455_ ), .ZN(\mycsreg/_0609_ ) );
NAND4_X1 \mycsreg/_1159_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0083_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0456_ ) );
NAND4_X1 \mycsreg/_1160_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0051_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0457_ ) );
NAND4_X1 \mycsreg/_1161_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0019_ ), .A3(\mycsreg/_0315_ ), .A4(\mycsreg/_0345_ ), .ZN(\mycsreg/_0458_ ) );
AND3_X1 \mycsreg/_1162_ ( .A1(\mycsreg/_0456_ ), .A2(\mycsreg/_0457_ ), .A3(\mycsreg/_0458_ ), .ZN(\mycsreg/_0459_ ) );
NAND4_X1 \mycsreg/_1163_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0115_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0460_ ) );
NAND3_X1 \mycsreg/_1164_ ( .A1(\mycsreg/_0459_ ), .A2(\mycsreg/_0330_ ), .A3(\mycsreg/_0460_ ), .ZN(\mycsreg/_0610_ ) );
AND4_X1 \mycsreg/_1165_ ( .A1(\mycsreg/_0052_ ), .A2(\mycsreg/_0277_ ), .A3(\mycsreg/_0344_ ), .A4(\mycsreg/_0283_ ), .ZN(\mycsreg/_0461_ ) );
AOI21_X1 \mycsreg/_1166_ ( .A(\mycsreg/_0461_ ), .B1(\mycsreg/_0275_ ), .B2(\mycsreg/_0297_ ), .ZN(\mycsreg/_0462_ ) );
NAND4_X1 \mycsreg/_1167_ ( .A1(\mycsreg/_0308_ ), .A2(\mycsreg/_0020_ ), .A3(\mycsreg/_0287_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0463_ ) );
NAND4_X1 \mycsreg/_1168_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0116_ ), .A3(\mycsreg/_0271_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0464_ ) );
NAND4_X1 \mycsreg/_1169_ ( .A1(\mycsreg/_0291_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0084_ ), .A4(\mycsreg/_0298_ ), .ZN(\mycsreg/_0465_ ) );
AND3_X1 \mycsreg/_1170_ ( .A1(\mycsreg/_0463_ ), .A2(\mycsreg/_0464_ ), .A3(\mycsreg/_0465_ ), .ZN(\mycsreg/_0466_ ) );
NAND2_X1 \mycsreg/_1171_ ( .A1(\mycsreg/_0462_ ), .A2(\mycsreg/_0466_ ), .ZN(\mycsreg/_0611_ ) );
NAND4_X1 \mycsreg/_1172_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0117_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0467_ ) );
NAND4_X1 \mycsreg/_1173_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0085_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0468_ ) );
NAND4_X1 \mycsreg/_1174_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0053_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0316_ ), .ZN(\mycsreg/_0469_ ) );
AND3_X1 \mycsreg/_1175_ ( .A1(\mycsreg/_0467_ ), .A2(\mycsreg/_0468_ ), .A3(\mycsreg/_0469_ ), .ZN(\mycsreg/_0470_ ) );
NAND4_X1 \mycsreg/_1176_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0021_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0471_ ) );
NAND3_X1 \mycsreg/_1177_ ( .A1(\mycsreg/_0470_ ), .A2(\mycsreg/_0330_ ), .A3(\mycsreg/_0471_ ), .ZN(\mycsreg/_0612_ ) );
NAND4_X1 \mycsreg/_1178_ ( .A1(\mycsreg/_0286_ ), .A2(\mycsreg/_0119_ ), .A3(\mycsreg/_0309_ ), .A4(\mycsreg/_0338_ ), .ZN(\mycsreg/_0472_ ) );
NAND4_X1 \mycsreg/_1179_ ( .A1(\mycsreg/_0312_ ), .A2(\mycsreg/_0296_ ), .A3(\mycsreg/_0087_ ), .A4(\mycsreg/_0292_ ), .ZN(\mycsreg/_0473_ ) );
NAND4_X1 \mycsreg/_1180_ ( .A1(\mycsreg/_0304_ ), .A2(\mycsreg/_0055_ ), .A3(\mycsreg/_0358_ ), .A4(\mycsreg/_0359_ ), .ZN(\mycsreg/_0474_ ) );
AND3_X1 \mycsreg/_1181_ ( .A1(\mycsreg/_0472_ ), .A2(\mycsreg/_0473_ ), .A3(\mycsreg/_0474_ ), .ZN(\mycsreg/_0475_ ) );
NAND4_X1 \mycsreg/_1182_ ( .A1(\mycsreg/_0301_ ), .A2(\mycsreg/_0023_ ), .A3(\mycsreg/_0302_ ), .A4(\mycsreg/_0322_ ), .ZN(\mycsreg/_0476_ ) );
NAND3_X1 \mycsreg/_1183_ ( .A1(\mycsreg/_0475_ ), .A2(\mycsreg/_0330_ ), .A3(\mycsreg/_0476_ ), .ZN(\mycsreg/_0614_ ) );
NAND4_X1 \mycsreg/_1184_ ( .A1(\mycsreg/_0295_ ), .A2(\mycsreg/_0120_ ), .A3(\mycsreg/_0272_ ), .A4(\mycsreg/_0299_ ), .ZN(\mycsreg/_0477_ ) );
NAND4_X1 \mycsreg/_1185_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0024_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0289_ ), .ZN(\mycsreg/_0478_ ) );
NAND4_X1 \mycsreg/_1186_ ( .A1(\mycsreg/_0305_ ), .A2(\mycsreg/_0313_ ), .A3(\mycsreg/_0088_ ), .A4(\mycsreg/_0310_ ), .ZN(\mycsreg/_0479_ ) );
NAND4_X1 \mycsreg/_1187_ ( .A1(\mycsreg/_0278_ ), .A2(\mycsreg/_0056_ ), .A3(\mycsreg/_0281_ ), .A4(\mycsreg/_0284_ ), .ZN(\mycsreg/_0480_ ) );
NAND4_X1 \mycsreg/_1188_ ( .A1(\mycsreg/_0477_ ), .A2(\mycsreg/_0478_ ), .A3(\mycsreg/_0479_ ), .A4(\mycsreg/_0480_ ), .ZN(\mycsreg/_0615_ ) );
MUX2_X1 \mycsreg/_1189_ ( .A(\mycsreg/_0636_ ), .B(\mycsreg/_0668_ ), .S(fanout_net_4 ), .Z(\mycsreg/_0481_ ) );
NOR2_X4 \mycsreg/_1190_ ( .A1(\mycsreg/_0631_ ), .A2(\mycsreg/_0630_ ), .ZN(\mycsreg/_0482_ ) );
INV_X1 \mycsreg/_1191_ ( .A(\mycsreg/_0633_ ), .ZN(\mycsreg/_0483_ ) );
NAND3_X2 \mycsreg/_1192_ ( .A1(\mycsreg/_0482_ ), .A2(\mycsreg/_0483_ ), .A3(\mycsreg/_0632_ ), .ZN(\mycsreg/_0484_ ) );
NOR2_X4 \mycsreg/_1193_ ( .A1(\mycsreg/_0629_ ), .A2(\mycsreg/_0628_ ), .ZN(\mycsreg/_0485_ ) );
INV_X2 \mycsreg/_1194_ ( .A(\mycsreg/_0485_ ), .ZN(\mycsreg/_0486_ ) );
INV_X1 \mycsreg/_1195_ ( .A(\mycsreg/_0627_ ), .ZN(\mycsreg/_0487_ ) );
NOR4_X2 \mycsreg/_1196_ ( .A1(\mycsreg/_0484_ ), .A2(\mycsreg/_0486_ ), .A3(\mycsreg/_0624_ ), .A4(\mycsreg/_0487_ ), .ZN(\mycsreg/_0488_ ) );
AND2_X1 \mycsreg/_1197_ ( .A1(\mycsreg/_0635_ ), .A2(\mycsreg/_0634_ ), .ZN(\mycsreg/_0489_ ) );
NOR2_X1 \mycsreg/_1198_ ( .A1(\mycsreg/_0626_ ), .A2(\mycsreg/_0625_ ), .ZN(\mycsreg/_0490_ ) );
AND3_X2 \mycsreg/_1199_ ( .A1(\mycsreg/_0488_ ), .A2(\mycsreg/_0489_ ), .A3(\mycsreg/_0490_ ), .ZN(\mycsreg/_0491_ ) );
OAI21_X2 \mycsreg/_1200_ ( .A(\mycsreg/_0675_ ), .B1(\mycsreg/_0491_ ), .B2(fanout_net_4 ), .ZN(\mycsreg/_0492_ ) );
NOR2_X4 \mycsreg/_1201_ ( .A1(\mycsreg/_0492_ ), .A2(\mycsreg/_0623_ ), .ZN(\mycsreg/_0493_ ) );
BUF_X4 \mycsreg/_1202_ ( .A(\mycsreg/_0493_ ), .Z(\mycsreg/_0494_ ) );
MUX2_X1 \mycsreg/_1203_ ( .A(\mycsreg/_0096_ ), .B(\mycsreg/_0481_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0128_ ) );
MUX2_X1 \mycsreg/_1204_ ( .A(\mycsreg/_0647_ ), .B(\mycsreg/_0669_ ), .S(fanout_net_4 ), .Z(\mycsreg/_0495_ ) );
MUX2_X1 \mycsreg/_1205_ ( .A(\mycsreg/_0107_ ), .B(\mycsreg/_0495_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0129_ ) );
MUX2_X1 \mycsreg/_1206_ ( .A(\mycsreg/_0658_ ), .B(\mycsreg/_0670_ ), .S(fanout_net_4 ), .Z(\mycsreg/_0496_ ) );
MUX2_X1 \mycsreg/_1207_ ( .A(\mycsreg/_0118_ ), .B(\mycsreg/_0496_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0130_ ) );
MUX2_X1 \mycsreg/_1208_ ( .A(\mycsreg/_0661_ ), .B(\mycsreg/_0671_ ), .S(fanout_net_4 ), .Z(\mycsreg/_0497_ ) );
MUX2_X1 \mycsreg/_1209_ ( .A(\mycsreg/_0121_ ), .B(\mycsreg/_0497_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0131_ ) );
MUX2_X1 \mycsreg/_1210_ ( .A(\mycsreg/_0662_ ), .B(\mycsreg/_0672_ ), .S(fanout_net_4 ), .Z(\mycsreg/_0498_ ) );
MUX2_X1 \mycsreg/_1211_ ( .A(\mycsreg/_0122_ ), .B(\mycsreg/_0498_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0132_ ) );
MUX2_X1 \mycsreg/_1212_ ( .A(\mycsreg/_0663_ ), .B(\mycsreg/_0673_ ), .S(fanout_net_4 ), .Z(\mycsreg/_0499_ ) );
MUX2_X1 \mycsreg/_1213_ ( .A(\mycsreg/_0123_ ), .B(\mycsreg/_0499_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0133_ ) );
INV_X1 \mycsreg/_1214_ ( .A(\mycsreg/_0482_ ), .ZN(\mycsreg/_0500_ ) );
OR3_X1 \mycsreg/_1215_ ( .A1(\mycsreg/_0500_ ), .A2(\mycsreg/_0633_ ), .A3(\mycsreg/_0632_ ), .ZN(\mycsreg/_0501_ ) );
NAND2_X1 \mycsreg/_1216_ ( .A1(\mycsreg/_0489_ ), .A2(\mycsreg/_0490_ ), .ZN(\mycsreg/_0502_ ) );
NOR2_X1 \mycsreg/_1217_ ( .A1(\mycsreg/_0501_ ), .A2(\mycsreg/_0502_ ), .ZN(\mycsreg/_0503_ ) );
INV_X1 \mycsreg/_1218_ ( .A(\mycsreg/_0675_ ), .ZN(\mycsreg/_0504_ ) );
NOR2_X1 \mycsreg/_1219_ ( .A1(\mycsreg/_0504_ ), .A2(\mycsreg/_0623_ ), .ZN(\mycsreg/_0505_ ) );
INV_X1 \mycsreg/_1220_ ( .A(\mycsreg/_0505_ ), .ZN(\mycsreg/_0506_ ) );
NOR4_X1 \mycsreg/_1221_ ( .A1(\mycsreg/_0506_ ), .A2(\mycsreg/_0486_ ), .A3(\mycsreg/_0624_ ), .A4(\mycsreg/_0627_ ), .ZN(\mycsreg/_0507_ ) );
NAND2_X1 \mycsreg/_1222_ ( .A1(\mycsreg/_0503_ ), .A2(\mycsreg/_0507_ ), .ZN(\mycsreg/_0508_ ) );
BUF_X4 \mycsreg/_1223_ ( .A(\mycsreg/_0508_ ), .Z(\mycsreg/_0509_ ) );
MUX2_X1 \mycsreg/_1224_ ( .A(\mycsreg/_0636_ ), .B(\mycsreg/_0000_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0134_ ) );
MUX2_X1 \mycsreg/_1225_ ( .A(\mycsreg/_0647_ ), .B(\mycsreg/_0011_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0135_ ) );
MUX2_X1 \mycsreg/_1226_ ( .A(\mycsreg/_0658_ ), .B(\mycsreg/_0022_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0136_ ) );
MUX2_X1 \mycsreg/_1227_ ( .A(\mycsreg/_0661_ ), .B(\mycsreg/_0025_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0137_ ) );
MUX2_X1 \mycsreg/_1228_ ( .A(\mycsreg/_0662_ ), .B(\mycsreg/_0026_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0138_ ) );
MUX2_X1 \mycsreg/_1229_ ( .A(\mycsreg/_0663_ ), .B(\mycsreg/_0027_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0139_ ) );
MUX2_X1 \mycsreg/_1230_ ( .A(\mycsreg/_0664_ ), .B(\mycsreg/_0028_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0140_ ) );
MUX2_X1 \mycsreg/_1231_ ( .A(\mycsreg/_0665_ ), .B(\mycsreg/_0029_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0141_ ) );
MUX2_X1 \mycsreg/_1232_ ( .A(\mycsreg/_0666_ ), .B(\mycsreg/_0030_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0142_ ) );
MUX2_X1 \mycsreg/_1233_ ( .A(\mycsreg/_0667_ ), .B(\mycsreg/_0031_ ), .S(\mycsreg/_0509_ ), .Z(\mycsreg/_0143_ ) );
BUF_X4 \mycsreg/_1234_ ( .A(\mycsreg/_0508_ ), .Z(\mycsreg/_0510_ ) );
MUX2_X1 \mycsreg/_1235_ ( .A(\mycsreg/_0637_ ), .B(\mycsreg/_0001_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0144_ ) );
MUX2_X1 \mycsreg/_1236_ ( .A(\mycsreg/_0638_ ), .B(\mycsreg/_0002_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0145_ ) );
MUX2_X1 \mycsreg/_1237_ ( .A(\mycsreg/_0639_ ), .B(\mycsreg/_0003_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0146_ ) );
MUX2_X1 \mycsreg/_1238_ ( .A(\mycsreg/_0640_ ), .B(\mycsreg/_0004_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0147_ ) );
MUX2_X1 \mycsreg/_1239_ ( .A(\mycsreg/_0641_ ), .B(\mycsreg/_0005_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0148_ ) );
MUX2_X1 \mycsreg/_1240_ ( .A(\mycsreg/_0642_ ), .B(\mycsreg/_0006_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0149_ ) );
MUX2_X1 \mycsreg/_1241_ ( .A(\mycsreg/_0643_ ), .B(\mycsreg/_0007_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0150_ ) );
MUX2_X1 \mycsreg/_1242_ ( .A(\mycsreg/_0644_ ), .B(\mycsreg/_0008_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0151_ ) );
MUX2_X1 \mycsreg/_1243_ ( .A(\mycsreg/_0645_ ), .B(\mycsreg/_0009_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0152_ ) );
MUX2_X1 \mycsreg/_1244_ ( .A(\mycsreg/_0646_ ), .B(\mycsreg/_0010_ ), .S(\mycsreg/_0510_ ), .Z(\mycsreg/_0153_ ) );
BUF_X4 \mycsreg/_1245_ ( .A(\mycsreg/_0508_ ), .Z(\mycsreg/_0511_ ) );
MUX2_X1 \mycsreg/_1246_ ( .A(\mycsreg/_0648_ ), .B(\mycsreg/_0012_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0154_ ) );
MUX2_X1 \mycsreg/_1247_ ( .A(\mycsreg/_0649_ ), .B(\mycsreg/_0013_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0155_ ) );
MUX2_X1 \mycsreg/_1248_ ( .A(\mycsreg/_0650_ ), .B(\mycsreg/_0014_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0156_ ) );
MUX2_X1 \mycsreg/_1249_ ( .A(\mycsreg/_0651_ ), .B(\mycsreg/_0015_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0157_ ) );
MUX2_X1 \mycsreg/_1250_ ( .A(\mycsreg/_0652_ ), .B(\mycsreg/_0016_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0158_ ) );
MUX2_X1 \mycsreg/_1251_ ( .A(\mycsreg/_0653_ ), .B(\mycsreg/_0017_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0159_ ) );
MUX2_X1 \mycsreg/_1252_ ( .A(\mycsreg/_0654_ ), .B(\mycsreg/_0018_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0160_ ) );
MUX2_X1 \mycsreg/_1253_ ( .A(\mycsreg/_0655_ ), .B(\mycsreg/_0019_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0161_ ) );
MUX2_X1 \mycsreg/_1254_ ( .A(\mycsreg/_0656_ ), .B(\mycsreg/_0020_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0162_ ) );
MUX2_X1 \mycsreg/_1255_ ( .A(\mycsreg/_0657_ ), .B(\mycsreg/_0021_ ), .S(\mycsreg/_0511_ ), .Z(\mycsreg/_0163_ ) );
MUX2_X1 \mycsreg/_1256_ ( .A(\mycsreg/_0659_ ), .B(\mycsreg/_0023_ ), .S(\mycsreg/_0508_ ), .Z(\mycsreg/_0164_ ) );
MUX2_X1 \mycsreg/_1257_ ( .A(\mycsreg/_0660_ ), .B(\mycsreg/_0024_ ), .S(\mycsreg/_0508_ ), .Z(\mycsreg/_0165_ ) );
INV_X1 \mycsreg/_1258_ ( .A(\mycsreg/_0628_ ), .ZN(\mycsreg/_0512_ ) );
NOR4_X1 \mycsreg/_1259_ ( .A1(\mycsreg/_0504_ ), .A2(\mycsreg/_0512_ ), .A3(\mycsreg/_0623_ ), .A4(\mycsreg/_0629_ ), .ZN(\mycsreg/_0513_ ) );
AND3_X1 \mycsreg/_1260_ ( .A1(\mycsreg/_0513_ ), .A2(\mycsreg/_0624_ ), .A3(\mycsreg/_0487_ ), .ZN(\mycsreg/_0514_ ) );
NAND2_X1 \mycsreg/_1261_ ( .A1(\mycsreg/_0503_ ), .A2(\mycsreg/_0514_ ), .ZN(\mycsreg/_0515_ ) );
BUF_X4 \mycsreg/_1262_ ( .A(\mycsreg/_0515_ ), .Z(\mycsreg/_0516_ ) );
MUX2_X1 \mycsreg/_1263_ ( .A(\mycsreg/_0636_ ), .B(\mycsreg/_0032_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0166_ ) );
MUX2_X1 \mycsreg/_1264_ ( .A(\mycsreg/_0647_ ), .B(\mycsreg/_0043_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0167_ ) );
MUX2_X1 \mycsreg/_1265_ ( .A(\mycsreg/_0658_ ), .B(\mycsreg/_0054_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0168_ ) );
MUX2_X1 \mycsreg/_1266_ ( .A(\mycsreg/_0661_ ), .B(\mycsreg/_0057_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0169_ ) );
MUX2_X1 \mycsreg/_1267_ ( .A(\mycsreg/_0662_ ), .B(\mycsreg/_0058_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0170_ ) );
MUX2_X1 \mycsreg/_1268_ ( .A(\mycsreg/_0663_ ), .B(\mycsreg/_0059_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0171_ ) );
MUX2_X1 \mycsreg/_1269_ ( .A(\mycsreg/_0664_ ), .B(\mycsreg/_0060_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0172_ ) );
MUX2_X1 \mycsreg/_1270_ ( .A(\mycsreg/_0665_ ), .B(\mycsreg/_0061_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0173_ ) );
MUX2_X1 \mycsreg/_1271_ ( .A(\mycsreg/_0666_ ), .B(\mycsreg/_0062_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0174_ ) );
MUX2_X1 \mycsreg/_1272_ ( .A(\mycsreg/_0667_ ), .B(\mycsreg/_0063_ ), .S(\mycsreg/_0516_ ), .Z(\mycsreg/_0175_ ) );
BUF_X4 \mycsreg/_1273_ ( .A(\mycsreg/_0515_ ), .Z(\mycsreg/_0517_ ) );
MUX2_X1 \mycsreg/_1274_ ( .A(\mycsreg/_0637_ ), .B(\mycsreg/_0033_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0176_ ) );
MUX2_X1 \mycsreg/_1275_ ( .A(\mycsreg/_0638_ ), .B(\mycsreg/_0034_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0177_ ) );
MUX2_X1 \mycsreg/_1276_ ( .A(\mycsreg/_0639_ ), .B(\mycsreg/_0035_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0178_ ) );
MUX2_X1 \mycsreg/_1277_ ( .A(\mycsreg/_0640_ ), .B(\mycsreg/_0036_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0179_ ) );
MUX2_X1 \mycsreg/_1278_ ( .A(\mycsreg/_0641_ ), .B(\mycsreg/_0037_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0180_ ) );
MUX2_X1 \mycsreg/_1279_ ( .A(\mycsreg/_0642_ ), .B(\mycsreg/_0038_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0181_ ) );
MUX2_X1 \mycsreg/_1280_ ( .A(\mycsreg/_0643_ ), .B(\mycsreg/_0039_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0182_ ) );
MUX2_X1 \mycsreg/_1281_ ( .A(\mycsreg/_0644_ ), .B(\mycsreg/_0040_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0183_ ) );
MUX2_X1 \mycsreg/_1282_ ( .A(\mycsreg/_0645_ ), .B(\mycsreg/_0041_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0184_ ) );
MUX2_X1 \mycsreg/_1283_ ( .A(\mycsreg/_0646_ ), .B(\mycsreg/_0042_ ), .S(\mycsreg/_0517_ ), .Z(\mycsreg/_0185_ ) );
BUF_X4 \mycsreg/_1284_ ( .A(\mycsreg/_0515_ ), .Z(\mycsreg/_0518_ ) );
MUX2_X1 \mycsreg/_1285_ ( .A(\mycsreg/_0648_ ), .B(\mycsreg/_0044_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0186_ ) );
MUX2_X1 \mycsreg/_1286_ ( .A(\mycsreg/_0649_ ), .B(\mycsreg/_0045_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0187_ ) );
MUX2_X1 \mycsreg/_1287_ ( .A(\mycsreg/_0650_ ), .B(\mycsreg/_0046_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0188_ ) );
MUX2_X1 \mycsreg/_1288_ ( .A(\mycsreg/_0651_ ), .B(\mycsreg/_0047_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0189_ ) );
MUX2_X1 \mycsreg/_1289_ ( .A(\mycsreg/_0652_ ), .B(\mycsreg/_0048_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0190_ ) );
MUX2_X1 \mycsreg/_1290_ ( .A(\mycsreg/_0653_ ), .B(\mycsreg/_0049_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0191_ ) );
MUX2_X1 \mycsreg/_1291_ ( .A(\mycsreg/_0654_ ), .B(\mycsreg/_0050_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0192_ ) );
MUX2_X1 \mycsreg/_1292_ ( .A(\mycsreg/_0655_ ), .B(\mycsreg/_0051_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0193_ ) );
MUX2_X1 \mycsreg/_1293_ ( .A(\mycsreg/_0656_ ), .B(\mycsreg/_0052_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0194_ ) );
MUX2_X1 \mycsreg/_1294_ ( .A(\mycsreg/_0657_ ), .B(\mycsreg/_0053_ ), .S(\mycsreg/_0518_ ), .Z(\mycsreg/_0195_ ) );
MUX2_X1 \mycsreg/_1295_ ( .A(\mycsreg/_0659_ ), .B(\mycsreg/_0055_ ), .S(\mycsreg/_0515_ ), .Z(\mycsreg/_0196_ ) );
MUX2_X1 \mycsreg/_1296_ ( .A(\mycsreg/_0660_ ), .B(\mycsreg/_0056_ ), .S(\mycsreg/_0515_ ), .Z(\mycsreg/_0197_ ) );
INV_X1 \mycsreg/_1297_ ( .A(\mycsreg/_0664_ ), .ZN(\mycsreg/_0519_ ) );
NOR2_X1 \mycsreg/_1298_ ( .A1(\mycsreg/_0519_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0520_ ) );
MUX2_X1 \mycsreg/_1299_ ( .A(\mycsreg/_0124_ ), .B(\mycsreg/_0520_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0198_ ) );
INV_X1 \mycsreg/_1300_ ( .A(\mycsreg/_0665_ ), .ZN(\mycsreg/_0521_ ) );
NOR2_X1 \mycsreg/_1301_ ( .A1(\mycsreg/_0521_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0522_ ) );
MUX2_X1 \mycsreg/_1302_ ( .A(\mycsreg/_0125_ ), .B(\mycsreg/_0522_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0199_ ) );
INV_X1 \mycsreg/_1303_ ( .A(\mycsreg/_0666_ ), .ZN(\mycsreg/_0523_ ) );
NOR2_X1 \mycsreg/_1304_ ( .A1(\mycsreg/_0523_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0524_ ) );
MUX2_X1 \mycsreg/_1305_ ( .A(\mycsreg/_0126_ ), .B(\mycsreg/_0524_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0200_ ) );
INV_X1 \mycsreg/_1306_ ( .A(\mycsreg/_0667_ ), .ZN(\mycsreg/_0525_ ) );
NOR2_X1 \mycsreg/_1307_ ( .A1(\mycsreg/_0525_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0526_ ) );
MUX2_X1 \mycsreg/_1308_ ( .A(\mycsreg/_0127_ ), .B(\mycsreg/_0526_ ), .S(\mycsreg/_0494_ ), .Z(\mycsreg/_0201_ ) );
INV_X1 \mycsreg/_1309_ ( .A(\mycsreg/_0637_ ), .ZN(\mycsreg/_0527_ ) );
NOR2_X1 \mycsreg/_1310_ ( .A1(\mycsreg/_0527_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0528_ ) );
BUF_X4 \mycsreg/_1311_ ( .A(\mycsreg/_0493_ ), .Z(\mycsreg/_0529_ ) );
MUX2_X1 \mycsreg/_1312_ ( .A(\mycsreg/_0097_ ), .B(\mycsreg/_0528_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0202_ ) );
INV_X1 \mycsreg/_1313_ ( .A(\mycsreg/_0638_ ), .ZN(\mycsreg/_0530_ ) );
NOR2_X1 \mycsreg/_1314_ ( .A1(\mycsreg/_0530_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0531_ ) );
MUX2_X1 \mycsreg/_1315_ ( .A(\mycsreg/_0098_ ), .B(\mycsreg/_0531_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0203_ ) );
INV_X1 \mycsreg/_1316_ ( .A(\mycsreg/_0639_ ), .ZN(\mycsreg/_0532_ ) );
NOR2_X1 \mycsreg/_1317_ ( .A1(\mycsreg/_0532_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0533_ ) );
MUX2_X1 \mycsreg/_1318_ ( .A(\mycsreg/_0099_ ), .B(\mycsreg/_0533_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0204_ ) );
INV_X1 \mycsreg/_1319_ ( .A(\mycsreg/_0640_ ), .ZN(\mycsreg/_0534_ ) );
NOR2_X1 \mycsreg/_1320_ ( .A1(\mycsreg/_0534_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0535_ ) );
MUX2_X1 \mycsreg/_1321_ ( .A(\mycsreg/_0100_ ), .B(\mycsreg/_0535_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0205_ ) );
INV_X1 \mycsreg/_1322_ ( .A(\mycsreg/_0641_ ), .ZN(\mycsreg/_0536_ ) );
NOR2_X1 \mycsreg/_1323_ ( .A1(\mycsreg/_0536_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0537_ ) );
MUX2_X1 \mycsreg/_1324_ ( .A(\mycsreg/_0101_ ), .B(\mycsreg/_0537_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0206_ ) );
INV_X1 \mycsreg/_1325_ ( .A(\mycsreg/_0642_ ), .ZN(\mycsreg/_0538_ ) );
NOR2_X1 \mycsreg/_1326_ ( .A1(\mycsreg/_0538_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0539_ ) );
MUX2_X1 \mycsreg/_1327_ ( .A(\mycsreg/_0102_ ), .B(\mycsreg/_0539_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0207_ ) );
INV_X1 \mycsreg/_1328_ ( .A(\mycsreg/_0643_ ), .ZN(\mycsreg/_0540_ ) );
NOR2_X1 \mycsreg/_1329_ ( .A1(\mycsreg/_0540_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0541_ ) );
MUX2_X1 \mycsreg/_1330_ ( .A(\mycsreg/_0103_ ), .B(\mycsreg/_0541_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0208_ ) );
INV_X1 \mycsreg/_1331_ ( .A(\mycsreg/_0644_ ), .ZN(\mycsreg/_0542_ ) );
NOR2_X1 \mycsreg/_1332_ ( .A1(\mycsreg/_0542_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0543_ ) );
MUX2_X1 \mycsreg/_1333_ ( .A(\mycsreg/_0104_ ), .B(\mycsreg/_0543_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0209_ ) );
INV_X1 \mycsreg/_1334_ ( .A(\mycsreg/_0645_ ), .ZN(\mycsreg/_0544_ ) );
NOR2_X1 \mycsreg/_1335_ ( .A1(\mycsreg/_0544_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0545_ ) );
MUX2_X1 \mycsreg/_1336_ ( .A(\mycsreg/_0105_ ), .B(\mycsreg/_0545_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0210_ ) );
INV_X1 \mycsreg/_1337_ ( .A(\mycsreg/_0646_ ), .ZN(\mycsreg/_0546_ ) );
NOR2_X1 \mycsreg/_1338_ ( .A1(\mycsreg/_0546_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0547_ ) );
MUX2_X1 \mycsreg/_1339_ ( .A(\mycsreg/_0106_ ), .B(\mycsreg/_0547_ ), .S(\mycsreg/_0529_ ), .Z(\mycsreg/_0211_ ) );
INV_X1 \mycsreg/_1340_ ( .A(\mycsreg/_0648_ ), .ZN(\mycsreg/_0548_ ) );
NOR2_X1 \mycsreg/_1341_ ( .A1(\mycsreg/_0548_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0549_ ) );
BUF_X4 \mycsreg/_1342_ ( .A(\mycsreg/_0493_ ), .Z(\mycsreg/_0550_ ) );
MUX2_X1 \mycsreg/_1343_ ( .A(\mycsreg/_0108_ ), .B(\mycsreg/_0549_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0212_ ) );
INV_X1 \mycsreg/_1344_ ( .A(\mycsreg/_0649_ ), .ZN(\mycsreg/_0551_ ) );
NOR2_X1 \mycsreg/_1345_ ( .A1(\mycsreg/_0551_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0552_ ) );
MUX2_X1 \mycsreg/_1346_ ( .A(\mycsreg/_0109_ ), .B(\mycsreg/_0552_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0213_ ) );
INV_X1 \mycsreg/_1347_ ( .A(\mycsreg/_0650_ ), .ZN(\mycsreg/_0553_ ) );
NOR2_X1 \mycsreg/_1348_ ( .A1(\mycsreg/_0553_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0554_ ) );
MUX2_X1 \mycsreg/_1349_ ( .A(\mycsreg/_0110_ ), .B(\mycsreg/_0554_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0214_ ) );
INV_X1 \mycsreg/_1350_ ( .A(\mycsreg/_0651_ ), .ZN(\mycsreg/_0555_ ) );
NOR2_X1 \mycsreg/_1351_ ( .A1(\mycsreg/_0555_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0556_ ) );
MUX2_X1 \mycsreg/_1352_ ( .A(\mycsreg/_0111_ ), .B(\mycsreg/_0556_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0215_ ) );
INV_X1 \mycsreg/_1353_ ( .A(\mycsreg/_0652_ ), .ZN(\mycsreg/_0557_ ) );
NOR2_X1 \mycsreg/_1354_ ( .A1(\mycsreg/_0557_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0558_ ) );
MUX2_X1 \mycsreg/_1355_ ( .A(\mycsreg/_0112_ ), .B(\mycsreg/_0558_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0216_ ) );
INV_X1 \mycsreg/_1356_ ( .A(\mycsreg/_0653_ ), .ZN(\mycsreg/_0559_ ) );
NOR2_X1 \mycsreg/_1357_ ( .A1(\mycsreg/_0559_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0560_ ) );
MUX2_X1 \mycsreg/_1358_ ( .A(\mycsreg/_0113_ ), .B(\mycsreg/_0560_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0217_ ) );
INV_X1 \mycsreg/_1359_ ( .A(\mycsreg/_0654_ ), .ZN(\mycsreg/_0561_ ) );
NOR2_X1 \mycsreg/_1360_ ( .A1(\mycsreg/_0561_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0562_ ) );
MUX2_X1 \mycsreg/_1361_ ( .A(\mycsreg/_0114_ ), .B(\mycsreg/_0562_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0218_ ) );
INV_X1 \mycsreg/_1362_ ( .A(\mycsreg/_0655_ ), .ZN(\mycsreg/_0563_ ) );
NOR2_X1 \mycsreg/_1363_ ( .A1(\mycsreg/_0563_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0564_ ) );
MUX2_X1 \mycsreg/_1364_ ( .A(\mycsreg/_0115_ ), .B(\mycsreg/_0564_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0219_ ) );
INV_X1 \mycsreg/_1365_ ( .A(\mycsreg/_0656_ ), .ZN(\mycsreg/_0565_ ) );
NOR2_X1 \mycsreg/_1366_ ( .A1(\mycsreg/_0565_ ), .A2(fanout_net_4 ), .ZN(\mycsreg/_0566_ ) );
MUX2_X1 \mycsreg/_1367_ ( .A(\mycsreg/_0116_ ), .B(\mycsreg/_0566_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0220_ ) );
INV_X1 \mycsreg/_1368_ ( .A(\mycsreg/_0657_ ), .ZN(\mycsreg/_0567_ ) );
NOR2_X1 \mycsreg/_1369_ ( .A1(\mycsreg/_0567_ ), .A2(\mycsreg/_0674_ ), .ZN(\mycsreg/_0568_ ) );
MUX2_X1 \mycsreg/_1370_ ( .A(\mycsreg/_0117_ ), .B(\mycsreg/_0568_ ), .S(\mycsreg/_0550_ ), .Z(\mycsreg/_0221_ ) );
INV_X1 \mycsreg/_1371_ ( .A(\mycsreg/_0659_ ), .ZN(\mycsreg/_0569_ ) );
NOR2_X1 \mycsreg/_1372_ ( .A1(\mycsreg/_0569_ ), .A2(\mycsreg/_0674_ ), .ZN(\mycsreg/_0570_ ) );
MUX2_X1 \mycsreg/_1373_ ( .A(\mycsreg/_0119_ ), .B(\mycsreg/_0570_ ), .S(\mycsreg/_0493_ ), .Z(\mycsreg/_0222_ ) );
INV_X1 \mycsreg/_1374_ ( .A(\mycsreg/_0660_ ), .ZN(\mycsreg/_0571_ ) );
NOR2_X1 \mycsreg/_1375_ ( .A1(\mycsreg/_0571_ ), .A2(\mycsreg/_0674_ ), .ZN(\mycsreg/_0572_ ) );
MUX2_X1 \mycsreg/_1376_ ( .A(\mycsreg/_0120_ ), .B(\mycsreg/_0572_ ), .S(\mycsreg/_0493_ ), .Z(\mycsreg/_0223_ ) );
AND4_X1 \mycsreg/_1377_ ( .A1(\mycsreg/_0624_ ), .A2(\mycsreg/_0505_ ), .A3(\mycsreg/_0487_ ), .A4(\mycsreg/_0485_ ), .ZN(\mycsreg/_0573_ ) );
NOR2_X1 \mycsreg/_1378_ ( .A1(\mycsreg/_0484_ ), .A2(\mycsreg/_0502_ ), .ZN(\mycsreg/_0574_ ) );
NAND2_X1 \mycsreg/_1379_ ( .A1(\mycsreg/_0573_ ), .A2(\mycsreg/_0574_ ), .ZN(\mycsreg/_0575_ ) );
BUF_X4 \mycsreg/_1380_ ( .A(\mycsreg/_0575_ ), .Z(\mycsreg/_0576_ ) );
MUX2_X1 \mycsreg/_1381_ ( .A(\mycsreg/_0636_ ), .B(\mycsreg/_0064_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0224_ ) );
MUX2_X1 \mycsreg/_1382_ ( .A(\mycsreg/_0647_ ), .B(\mycsreg/_0075_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0225_ ) );
MUX2_X1 \mycsreg/_1383_ ( .A(\mycsreg/_0658_ ), .B(\mycsreg/_0086_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0226_ ) );
MUX2_X1 \mycsreg/_1384_ ( .A(\mycsreg/_0661_ ), .B(\mycsreg/_0089_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0227_ ) );
MUX2_X1 \mycsreg/_1385_ ( .A(\mycsreg/_0662_ ), .B(\mycsreg/_0090_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0228_ ) );
MUX2_X1 \mycsreg/_1386_ ( .A(\mycsreg/_0663_ ), .B(\mycsreg/_0091_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0229_ ) );
MUX2_X1 \mycsreg/_1387_ ( .A(\mycsreg/_0664_ ), .B(\mycsreg/_0092_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0230_ ) );
MUX2_X1 \mycsreg/_1388_ ( .A(\mycsreg/_0665_ ), .B(\mycsreg/_0093_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0231_ ) );
MUX2_X1 \mycsreg/_1389_ ( .A(\mycsreg/_0666_ ), .B(\mycsreg/_0094_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0232_ ) );
MUX2_X1 \mycsreg/_1390_ ( .A(\mycsreg/_0667_ ), .B(\mycsreg/_0095_ ), .S(\mycsreg/_0576_ ), .Z(\mycsreg/_0233_ ) );
BUF_X4 \mycsreg/_1391_ ( .A(\mycsreg/_0575_ ), .Z(\mycsreg/_0577_ ) );
MUX2_X1 \mycsreg/_1392_ ( .A(\mycsreg/_0637_ ), .B(\mycsreg/_0065_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0234_ ) );
MUX2_X1 \mycsreg/_1393_ ( .A(\mycsreg/_0638_ ), .B(\mycsreg/_0066_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0235_ ) );
MUX2_X1 \mycsreg/_1394_ ( .A(\mycsreg/_0639_ ), .B(\mycsreg/_0067_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0236_ ) );
MUX2_X1 \mycsreg/_1395_ ( .A(\mycsreg/_0640_ ), .B(\mycsreg/_0068_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0237_ ) );
MUX2_X1 \mycsreg/_1396_ ( .A(\mycsreg/_0641_ ), .B(\mycsreg/_0069_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0238_ ) );
MUX2_X1 \mycsreg/_1397_ ( .A(\mycsreg/_0642_ ), .B(\mycsreg/_0070_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0239_ ) );
MUX2_X1 \mycsreg/_1398_ ( .A(\mycsreg/_0643_ ), .B(\mycsreg/_0071_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0240_ ) );
MUX2_X1 \mycsreg/_1399_ ( .A(\mycsreg/_0644_ ), .B(\mycsreg/_0072_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0241_ ) );
MUX2_X1 \mycsreg/_1400_ ( .A(\mycsreg/_0645_ ), .B(\mycsreg/_0073_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0242_ ) );
MUX2_X1 \mycsreg/_1401_ ( .A(\mycsreg/_0646_ ), .B(\mycsreg/_0074_ ), .S(\mycsreg/_0577_ ), .Z(\mycsreg/_0243_ ) );
BUF_X4 \mycsreg/_1402_ ( .A(\mycsreg/_0575_ ), .Z(\mycsreg/_0578_ ) );
MUX2_X1 \mycsreg/_1403_ ( .A(\mycsreg/_0648_ ), .B(\mycsreg/_0076_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0244_ ) );
MUX2_X1 \mycsreg/_1404_ ( .A(\mycsreg/_0649_ ), .B(\mycsreg/_0077_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0245_ ) );
MUX2_X1 \mycsreg/_1405_ ( .A(\mycsreg/_0650_ ), .B(\mycsreg/_0078_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0246_ ) );
MUX2_X1 \mycsreg/_1406_ ( .A(\mycsreg/_0651_ ), .B(\mycsreg/_0079_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0247_ ) );
MUX2_X1 \mycsreg/_1407_ ( .A(\mycsreg/_0652_ ), .B(\mycsreg/_0080_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0248_ ) );
MUX2_X1 \mycsreg/_1408_ ( .A(\mycsreg/_0653_ ), .B(\mycsreg/_0081_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0249_ ) );
MUX2_X1 \mycsreg/_1409_ ( .A(\mycsreg/_0654_ ), .B(\mycsreg/_0082_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0250_ ) );
MUX2_X1 \mycsreg/_1410_ ( .A(\mycsreg/_0655_ ), .B(\mycsreg/_0083_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0251_ ) );
MUX2_X1 \mycsreg/_1411_ ( .A(\mycsreg/_0656_ ), .B(\mycsreg/_0084_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0252_ ) );
MUX2_X1 \mycsreg/_1412_ ( .A(\mycsreg/_0657_ ), .B(\mycsreg/_0085_ ), .S(\mycsreg/_0578_ ), .Z(\mycsreg/_0253_ ) );
MUX2_X1 \mycsreg/_1413_ ( .A(\mycsreg/_0659_ ), .B(\mycsreg/_0087_ ), .S(\mycsreg/_0575_ ), .Z(\mycsreg/_0254_ ) );
MUX2_X1 \mycsreg/_1414_ ( .A(\mycsreg/_0660_ ), .B(\mycsreg/_0088_ ), .S(\mycsreg/_0575_ ), .Z(\mycsreg/_0255_ ) );
DFF_X1 \mycsreg/_1415_ ( .D(\mycsreg/_0804_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][0] ), .QN(\mycsreg/_0803_ ) );
DFF_X1 \mycsreg/_1416_ ( .D(\mycsreg/_0805_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][1] ), .QN(\mycsreg/_0802_ ) );
DFF_X1 \mycsreg/_1417_ ( .D(\mycsreg/_0806_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][2] ), .QN(\mycsreg/_0801_ ) );
DFF_X1 \mycsreg/_1418_ ( .D(\mycsreg/_0807_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][3] ), .QN(\mycsreg/_0800_ ) );
DFF_X1 \mycsreg/_1419_ ( .D(\mycsreg/_0808_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][4] ), .QN(\mycsreg/_0799_ ) );
DFF_X1 \mycsreg/_1420_ ( .D(\mycsreg/_0809_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][5] ), .QN(\mycsreg/_0798_ ) );
DFF_X1 \mycsreg/_1421_ ( .D(\mycsreg/_0810_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][0] ), .QN(\mycsreg/_0797_ ) );
DFF_X1 \mycsreg/_1422_ ( .D(\mycsreg/_0811_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][1] ), .QN(\mycsreg/_0796_ ) );
DFF_X1 \mycsreg/_1423_ ( .D(\mycsreg/_0812_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][2] ), .QN(\mycsreg/_0795_ ) );
DFF_X1 \mycsreg/_1424_ ( .D(\mycsreg/_0813_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][3] ), .QN(\mycsreg/_0794_ ) );
DFF_X1 \mycsreg/_1425_ ( .D(\mycsreg/_0814_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][4] ), .QN(\mycsreg/_0793_ ) );
DFF_X1 \mycsreg/_1426_ ( .D(\mycsreg/_0815_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][5] ), .QN(\mycsreg/_0792_ ) );
DFF_X1 \mycsreg/_1427_ ( .D(\mycsreg/_0816_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][6] ), .QN(\mycsreg/_0791_ ) );
DFF_X1 \mycsreg/_1428_ ( .D(\mycsreg/_0817_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][7] ), .QN(\mycsreg/_0790_ ) );
DFF_X1 \mycsreg/_1429_ ( .D(\mycsreg/_0818_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][8] ), .QN(\mycsreg/_0789_ ) );
DFF_X1 \mycsreg/_1430_ ( .D(\mycsreg/_0819_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][9] ), .QN(\mycsreg/_0788_ ) );
DFF_X1 \mycsreg/_1431_ ( .D(\mycsreg/_0820_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][10] ), .QN(\mycsreg/_0787_ ) );
DFF_X1 \mycsreg/_1432_ ( .D(\mycsreg/_0821_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][11] ), .QN(\mycsreg/_0786_ ) );
DFF_X1 \mycsreg/_1433_ ( .D(\mycsreg/_0822_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][12] ), .QN(\mycsreg/_0785_ ) );
DFF_X1 \mycsreg/_1434_ ( .D(\mycsreg/_0823_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][13] ), .QN(\mycsreg/_0784_ ) );
DFF_X1 \mycsreg/_1435_ ( .D(\mycsreg/_0824_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][14] ), .QN(\mycsreg/_0783_ ) );
DFF_X1 \mycsreg/_1436_ ( .D(\mycsreg/_0825_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][15] ), .QN(\mycsreg/_0782_ ) );
DFF_X1 \mycsreg/_1437_ ( .D(\mycsreg/_0826_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][16] ), .QN(\mycsreg/_0781_ ) );
DFF_X1 \mycsreg/_1438_ ( .D(\mycsreg/_0827_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][17] ), .QN(\mycsreg/_0780_ ) );
DFF_X1 \mycsreg/_1439_ ( .D(\mycsreg/_0828_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][18] ), .QN(\mycsreg/_0779_ ) );
DFF_X1 \mycsreg/_1440_ ( .D(\mycsreg/_0829_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][19] ), .QN(\mycsreg/_0778_ ) );
DFF_X1 \mycsreg/_1441_ ( .D(\mycsreg/_0830_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][20] ), .QN(\mycsreg/_0777_ ) );
DFF_X1 \mycsreg/_1442_ ( .D(\mycsreg/_0831_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][21] ), .QN(\mycsreg/_0776_ ) );
DFF_X1 \mycsreg/_1443_ ( .D(\mycsreg/_0832_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][22] ), .QN(\mycsreg/_0775_ ) );
DFF_X1 \mycsreg/_1444_ ( .D(\mycsreg/_0833_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][23] ), .QN(\mycsreg/_0774_ ) );
DFF_X1 \mycsreg/_1445_ ( .D(\mycsreg/_0834_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][24] ), .QN(\mycsreg/_0773_ ) );
DFF_X1 \mycsreg/_1446_ ( .D(\mycsreg/_0835_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][25] ), .QN(\mycsreg/_0772_ ) );
DFF_X1 \mycsreg/_1447_ ( .D(\mycsreg/_0836_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][26] ), .QN(\mycsreg/_0771_ ) );
DFF_X1 \mycsreg/_1448_ ( .D(\mycsreg/_0837_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][27] ), .QN(\mycsreg/_0770_ ) );
DFF_X1 \mycsreg/_1449_ ( .D(\mycsreg/_0838_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][28] ), .QN(\mycsreg/_0769_ ) );
DFF_X1 \mycsreg/_1450_ ( .D(\mycsreg/_0839_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][29] ), .QN(\mycsreg/_0768_ ) );
DFF_X1 \mycsreg/_1451_ ( .D(\mycsreg/_0840_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][30] ), .QN(\mycsreg/_0767_ ) );
DFF_X1 \mycsreg/_1452_ ( .D(\mycsreg/_0841_ ), .CK(clock ), .Q(\mycsreg/CSReg[0][31] ), .QN(\mycsreg/_0766_ ) );
DFF_X1 \mycsreg/_1453_ ( .D(\mycsreg/_0842_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][0] ), .QN(\mycsreg/_0765_ ) );
DFF_X1 \mycsreg/_1454_ ( .D(\mycsreg/_0843_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][1] ), .QN(\mycsreg/_0764_ ) );
DFF_X1 \mycsreg/_1455_ ( .D(\mycsreg/_0844_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][2] ), .QN(\mycsreg/_0763_ ) );
DFF_X1 \mycsreg/_1456_ ( .D(\mycsreg/_0845_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][3] ), .QN(\mycsreg/_0762_ ) );
DFF_X1 \mycsreg/_1457_ ( .D(\mycsreg/_0846_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][4] ), .QN(\mycsreg/_0761_ ) );
DFF_X1 \mycsreg/_1458_ ( .D(\mycsreg/_0847_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][5] ), .QN(\mycsreg/_0760_ ) );
DFF_X1 \mycsreg/_1459_ ( .D(\mycsreg/_0848_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][6] ), .QN(\mycsreg/_0759_ ) );
DFF_X1 \mycsreg/_1460_ ( .D(\mycsreg/_0849_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][7] ), .QN(\mycsreg/_0758_ ) );
DFF_X1 \mycsreg/_1461_ ( .D(\mycsreg/_0850_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][8] ), .QN(\mycsreg/_0757_ ) );
DFF_X1 \mycsreg/_1462_ ( .D(\mycsreg/_0851_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][9] ), .QN(\mycsreg/_0756_ ) );
DFF_X1 \mycsreg/_1463_ ( .D(\mycsreg/_0852_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][10] ), .QN(\mycsreg/_0755_ ) );
DFF_X1 \mycsreg/_1464_ ( .D(\mycsreg/_0853_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][11] ), .QN(\mycsreg/_0754_ ) );
DFF_X1 \mycsreg/_1465_ ( .D(\mycsreg/_0854_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][12] ), .QN(\mycsreg/_0753_ ) );
DFF_X1 \mycsreg/_1466_ ( .D(\mycsreg/_0855_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][13] ), .QN(\mycsreg/_0752_ ) );
DFF_X1 \mycsreg/_1467_ ( .D(\mycsreg/_0856_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][14] ), .QN(\mycsreg/_0751_ ) );
DFF_X1 \mycsreg/_1468_ ( .D(\mycsreg/_0857_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][15] ), .QN(\mycsreg/_0750_ ) );
DFF_X1 \mycsreg/_1469_ ( .D(\mycsreg/_0858_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][16] ), .QN(\mycsreg/_0749_ ) );
DFF_X1 \mycsreg/_1470_ ( .D(\mycsreg/_0859_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][17] ), .QN(\mycsreg/_0748_ ) );
DFF_X1 \mycsreg/_1471_ ( .D(\mycsreg/_0860_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][18] ), .QN(\mycsreg/_0747_ ) );
DFF_X1 \mycsreg/_1472_ ( .D(\mycsreg/_0861_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][19] ), .QN(\mycsreg/_0746_ ) );
DFF_X1 \mycsreg/_1473_ ( .D(\mycsreg/_0862_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][20] ), .QN(\mycsreg/_0745_ ) );
DFF_X1 \mycsreg/_1474_ ( .D(\mycsreg/_0863_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][21] ), .QN(\mycsreg/_0744_ ) );
DFF_X1 \mycsreg/_1475_ ( .D(\mycsreg/_0864_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][22] ), .QN(\mycsreg/_0743_ ) );
DFF_X1 \mycsreg/_1476_ ( .D(\mycsreg/_0865_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][23] ), .QN(\mycsreg/_0742_ ) );
DFF_X1 \mycsreg/_1477_ ( .D(\mycsreg/_0866_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][24] ), .QN(\mycsreg/_0741_ ) );
DFF_X1 \mycsreg/_1478_ ( .D(\mycsreg/_0867_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][25] ), .QN(\mycsreg/_0740_ ) );
DFF_X1 \mycsreg/_1479_ ( .D(\mycsreg/_0868_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][26] ), .QN(\mycsreg/_0739_ ) );
DFF_X1 \mycsreg/_1480_ ( .D(\mycsreg/_0869_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][27] ), .QN(\mycsreg/_0738_ ) );
DFF_X1 \mycsreg/_1481_ ( .D(\mycsreg/_0870_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][28] ), .QN(\mycsreg/_0737_ ) );
DFF_X1 \mycsreg/_1482_ ( .D(\mycsreg/_0871_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][29] ), .QN(\mycsreg/_0736_ ) );
DFF_X1 \mycsreg/_1483_ ( .D(\mycsreg/_0872_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][30] ), .QN(\mycsreg/_0735_ ) );
DFF_X1 \mycsreg/_1484_ ( .D(\mycsreg/_0873_ ), .CK(clock ), .Q(\mycsreg/CSReg[1][31] ), .QN(\mycsreg/_0734_ ) );
DFF_X1 \mycsreg/_1485_ ( .D(\mycsreg/_0874_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][6] ), .QN(\mycsreg/_0733_ ) );
DFF_X1 \mycsreg/_1486_ ( .D(\mycsreg/_0875_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][7] ), .QN(\mycsreg/_0732_ ) );
DFF_X1 \mycsreg/_1487_ ( .D(\mycsreg/_0876_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][8] ), .QN(\mycsreg/_0731_ ) );
DFF_X1 \mycsreg/_1488_ ( .D(\mycsreg/_0877_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][9] ), .QN(\mycsreg/_0730_ ) );
DFF_X1 \mycsreg/_1489_ ( .D(\mycsreg/_0878_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][10] ), .QN(\mycsreg/_0729_ ) );
DFF_X1 \mycsreg/_1490_ ( .D(\mycsreg/_0879_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][11] ), .QN(\mycsreg/_0728_ ) );
DFF_X1 \mycsreg/_1491_ ( .D(\mycsreg/_0880_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][12] ), .QN(\mycsreg/_0727_ ) );
DFF_X1 \mycsreg/_1492_ ( .D(\mycsreg/_0881_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][13] ), .QN(\mycsreg/_0726_ ) );
DFF_X1 \mycsreg/_1493_ ( .D(\mycsreg/_0882_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][14] ), .QN(\mycsreg/_0725_ ) );
DFF_X1 \mycsreg/_1494_ ( .D(\mycsreg/_0883_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][15] ), .QN(\mycsreg/_0724_ ) );
DFF_X1 \mycsreg/_1495_ ( .D(\mycsreg/_0884_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][16] ), .QN(\mycsreg/_0723_ ) );
DFF_X1 \mycsreg/_1496_ ( .D(\mycsreg/_0885_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][17] ), .QN(\mycsreg/_0722_ ) );
DFF_X1 \mycsreg/_1497_ ( .D(\mycsreg/_0886_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][18] ), .QN(\mycsreg/_0721_ ) );
DFF_X1 \mycsreg/_1498_ ( .D(\mycsreg/_0887_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][19] ), .QN(\mycsreg/_0720_ ) );
DFF_X1 \mycsreg/_1499_ ( .D(\mycsreg/_0888_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][20] ), .QN(\mycsreg/_0719_ ) );
DFF_X1 \mycsreg/_1500_ ( .D(\mycsreg/_0889_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][21] ), .QN(\mycsreg/_0718_ ) );
DFF_X1 \mycsreg/_1501_ ( .D(\mycsreg/_0890_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][22] ), .QN(\mycsreg/_0717_ ) );
DFF_X1 \mycsreg/_1502_ ( .D(\mycsreg/_0891_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][23] ), .QN(\mycsreg/_0716_ ) );
DFF_X1 \mycsreg/_1503_ ( .D(\mycsreg/_0892_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][24] ), .QN(\mycsreg/_0715_ ) );
DFF_X1 \mycsreg/_1504_ ( .D(\mycsreg/_0893_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][25] ), .QN(\mycsreg/_0714_ ) );
DFF_X1 \mycsreg/_1505_ ( .D(\mycsreg/_0894_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][26] ), .QN(\mycsreg/_0713_ ) );
DFF_X1 \mycsreg/_1506_ ( .D(\mycsreg/_0895_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][27] ), .QN(\mycsreg/_0712_ ) );
DFF_X1 \mycsreg/_1507_ ( .D(\mycsreg/_0896_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][28] ), .QN(\mycsreg/_0711_ ) );
DFF_X1 \mycsreg/_1508_ ( .D(\mycsreg/_0897_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][29] ), .QN(\mycsreg/_0710_ ) );
DFF_X1 \mycsreg/_1509_ ( .D(\mycsreg/_0898_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][30] ), .QN(\mycsreg/_0709_ ) );
DFF_X1 \mycsreg/_1510_ ( .D(\mycsreg/_0899_ ), .CK(clock ), .Q(\mycsreg/CSReg[3][31] ), .QN(\mycsreg/_0708_ ) );
DFF_X1 \mycsreg/_1511_ ( .D(\mycsreg/_0900_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][0] ), .QN(\mycsreg/_0707_ ) );
DFF_X1 \mycsreg/_1512_ ( .D(\mycsreg/_0901_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][1] ), .QN(\mycsreg/_0706_ ) );
DFF_X1 \mycsreg/_1513_ ( .D(\mycsreg/_0902_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][2] ), .QN(\mycsreg/_0705_ ) );
DFF_X1 \mycsreg/_1514_ ( .D(\mycsreg/_0903_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][3] ), .QN(\mycsreg/_0704_ ) );
DFF_X1 \mycsreg/_1515_ ( .D(\mycsreg/_0904_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][4] ), .QN(\mycsreg/_0703_ ) );
DFF_X1 \mycsreg/_1516_ ( .D(\mycsreg/_0905_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][5] ), .QN(\mycsreg/_0702_ ) );
DFF_X1 \mycsreg/_1517_ ( .D(\mycsreg/_0906_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][6] ), .QN(\mycsreg/_0701_ ) );
DFF_X1 \mycsreg/_1518_ ( .D(\mycsreg/_0907_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][7] ), .QN(\mycsreg/_0700_ ) );
DFF_X1 \mycsreg/_1519_ ( .D(\mycsreg/_0908_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][8] ), .QN(\mycsreg/_0699_ ) );
DFF_X1 \mycsreg/_1520_ ( .D(\mycsreg/_0909_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][9] ), .QN(\mycsreg/_0698_ ) );
DFF_X1 \mycsreg/_1521_ ( .D(\mycsreg/_0910_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][10] ), .QN(\mycsreg/_0697_ ) );
DFF_X1 \mycsreg/_1522_ ( .D(\mycsreg/_0911_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][11] ), .QN(\mycsreg/_0696_ ) );
DFF_X1 \mycsreg/_1523_ ( .D(\mycsreg/_0912_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][12] ), .QN(\mycsreg/_0695_ ) );
DFF_X1 \mycsreg/_1524_ ( .D(\mycsreg/_0913_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][13] ), .QN(\mycsreg/_0694_ ) );
DFF_X1 \mycsreg/_1525_ ( .D(\mycsreg/_0914_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][14] ), .QN(\mycsreg/_0693_ ) );
DFF_X1 \mycsreg/_1526_ ( .D(\mycsreg/_0915_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][15] ), .QN(\mycsreg/_0692_ ) );
DFF_X1 \mycsreg/_1527_ ( .D(\mycsreg/_0916_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][16] ), .QN(\mycsreg/_0691_ ) );
DFF_X1 \mycsreg/_1528_ ( .D(\mycsreg/_0917_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][17] ), .QN(\mycsreg/_0690_ ) );
DFF_X1 \mycsreg/_1529_ ( .D(\mycsreg/_0918_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][18] ), .QN(\mycsreg/_0689_ ) );
DFF_X1 \mycsreg/_1530_ ( .D(\mycsreg/_0919_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][19] ), .QN(\mycsreg/_0688_ ) );
DFF_X1 \mycsreg/_1531_ ( .D(\mycsreg/_0920_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][20] ), .QN(\mycsreg/_0687_ ) );
DFF_X1 \mycsreg/_1532_ ( .D(\mycsreg/_0921_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][21] ), .QN(\mycsreg/_0686_ ) );
DFF_X1 \mycsreg/_1533_ ( .D(\mycsreg/_0922_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][22] ), .QN(\mycsreg/_0685_ ) );
DFF_X1 \mycsreg/_1534_ ( .D(\mycsreg/_0923_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][23] ), .QN(\mycsreg/_0684_ ) );
DFF_X1 \mycsreg/_1535_ ( .D(\mycsreg/_0924_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][24] ), .QN(\mycsreg/_0683_ ) );
DFF_X1 \mycsreg/_1536_ ( .D(\mycsreg/_0925_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][25] ), .QN(\mycsreg/_0682_ ) );
DFF_X1 \mycsreg/_1537_ ( .D(\mycsreg/_0926_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][26] ), .QN(\mycsreg/_0681_ ) );
DFF_X1 \mycsreg/_1538_ ( .D(\mycsreg/_0927_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][27] ), .QN(\mycsreg/_0680_ ) );
DFF_X1 \mycsreg/_1539_ ( .D(\mycsreg/_0928_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][28] ), .QN(\mycsreg/_0679_ ) );
DFF_X1 \mycsreg/_1540_ ( .D(\mycsreg/_0929_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][29] ), .QN(\mycsreg/_0678_ ) );
DFF_X1 \mycsreg/_1541_ ( .D(\mycsreg/_0930_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][30] ), .QN(\mycsreg/_0677_ ) );
DFF_X1 \mycsreg/_1542_ ( .D(\mycsreg/_0931_ ), .CK(clock ), .Q(\mycsreg/CSReg[2][31] ), .QN(\mycsreg/_0676_ ) );
BUF_X1 \mycsreg/_1543_ ( .A(\LS_WB_wen_csreg [7] ), .Z(\mycsreg/_0675_ ) );
BUF_X1 \mycsreg/_1544_ ( .A(reset ), .Z(\mycsreg/_0623_ ) );
BUF_X1 \mycsreg/_1545_ ( .A(\LS_WB_waddr_csreg [0] ), .Z(\mycsreg/_0624_ ) );
BUF_X1 \mycsreg/_1546_ ( .A(\LS_WB_waddr_csreg [1] ), .Z(\mycsreg/_0627_ ) );
BUF_X1 \mycsreg/_1547_ ( .A(\LS_WB_waddr_csreg [3] ), .Z(\mycsreg/_0629_ ) );
BUF_X1 \mycsreg/_1548_ ( .A(\LS_WB_waddr_csreg [2] ), .Z(\mycsreg/_0628_ ) );
BUF_X1 \mycsreg/_1549_ ( .A(\LS_WB_waddr_csreg [5] ), .Z(\mycsreg/_0631_ ) );
BUF_X1 \mycsreg/_1550_ ( .A(\LS_WB_waddr_csreg [4] ), .Z(\mycsreg/_0630_ ) );
BUF_X1 \mycsreg/_1551_ ( .A(\LS_WB_waddr_csreg [7] ), .Z(\mycsreg/_0633_ ) );
BUF_X1 \mycsreg/_1552_ ( .A(\LS_WB_waddr_csreg [6] ), .Z(\mycsreg/_0632_ ) );
BUF_X1 \mycsreg/_1553_ ( .A(\LS_WB_waddr_csreg [9] ), .Z(\mycsreg/_0635_ ) );
BUF_X1 \mycsreg/_1554_ ( .A(\LS_WB_waddr_csreg [8] ), .Z(\mycsreg/_0634_ ) );
BUF_X1 \mycsreg/_1555_ ( .A(\LS_WB_waddr_csreg [11] ), .Z(\mycsreg/_0626_ ) );
BUF_X1 \mycsreg/_1556_ ( .A(\LS_WB_waddr_csreg [10] ), .Z(\mycsreg/_0625_ ) );
BUF_X1 \mycsreg/_1557_ ( .A(\LS_WB_wen_csreg [6] ), .Z(\mycsreg/_0674_ ) );
BUF_X1 \mycsreg/_1558_ ( .A(\ID_EX_csr [9] ), .Z(\mycsreg/_0590_ ) );
BUF_X1 \mycsreg/_1559_ ( .A(\ID_EX_csr [8] ), .Z(\mycsreg/_0589_ ) );
BUF_X1 \mycsreg/_1560_ ( .A(\ID_EX_csr [11] ), .Z(\mycsreg/_0581_ ) );
BUF_X1 \mycsreg/_1561_ ( .A(\ID_EX_csr [10] ), .Z(\mycsreg/_0580_ ) );
BUF_X1 \mycsreg/_1562_ ( .A(\ID_EX_csr [7] ), .Z(\mycsreg/_0588_ ) );
BUF_X1 \mycsreg/_1563_ ( .A(\ID_EX_csr [6] ), .Z(\mycsreg/_0587_ ) );
BUF_X1 \mycsreg/_1564_ ( .A(\ID_EX_csr [5] ), .Z(\mycsreg/_0586_ ) );
BUF_X1 \mycsreg/_1565_ ( .A(\ID_EX_csr [4] ), .Z(\mycsreg/_0585_ ) );
BUF_X1 \mycsreg/_1566_ ( .A(\ID_EX_csr [3] ), .Z(\mycsreg/_0584_ ) );
BUF_X1 \mycsreg/_1567_ ( .A(\ID_EX_csr [2] ), .Z(\mycsreg/_0583_ ) );
BUF_X1 \mycsreg/_1568_ ( .A(\ID_EX_csr [1] ), .Z(\mycsreg/_0582_ ) );
BUF_X1 \mycsreg/_1569_ ( .A(\ID_EX_csr [0] ), .Z(\mycsreg/_0579_ ) );
BUF_X1 \mycsreg/_1570_ ( .A(\mycsreg/CSReg[3][0] ), .Z(\mycsreg/_0096_ ) );
BUF_X1 \mycsreg/_1571_ ( .A(\mycsreg/CSReg[2][0] ), .Z(\mycsreg/_0064_ ) );
BUF_X1 \mycsreg/_1572_ ( .A(\mycsreg/CSReg[1][0] ), .Z(\mycsreg/_0032_ ) );
BUF_X1 \mycsreg/_1573_ ( .A(\mycsreg/CSReg[0][0] ), .Z(\mycsreg/_0000_ ) );
BUF_X1 \mycsreg/_1574_ ( .A(\mycsreg/_0591_ ), .Z(\srccs_raw [0] ) );
BUF_X1 \mycsreg/_1575_ ( .A(\mycsreg/CSReg[3][1] ), .Z(\mycsreg/_0107_ ) );
BUF_X1 \mycsreg/_1576_ ( .A(\mycsreg/CSReg[2][1] ), .Z(\mycsreg/_0075_ ) );
BUF_X1 \mycsreg/_1577_ ( .A(\mycsreg/CSReg[1][1] ), .Z(\mycsreg/_0043_ ) );
BUF_X1 \mycsreg/_1578_ ( .A(\mycsreg/CSReg[0][1] ), .Z(\mycsreg/_0011_ ) );
BUF_X1 \mycsreg/_1579_ ( .A(\mycsreg/_0602_ ), .Z(\srccs_raw [1] ) );
BUF_X1 \mycsreg/_1580_ ( .A(\mycsreg/CSReg[3][2] ), .Z(\mycsreg/_0118_ ) );
BUF_X1 \mycsreg/_1581_ ( .A(\mycsreg/CSReg[2][2] ), .Z(\mycsreg/_0086_ ) );
BUF_X1 \mycsreg/_1582_ ( .A(\mycsreg/CSReg[1][2] ), .Z(\mycsreg/_0054_ ) );
BUF_X1 \mycsreg/_1583_ ( .A(\mycsreg/CSReg[0][2] ), .Z(\mycsreg/_0022_ ) );
BUF_X1 \mycsreg/_1584_ ( .A(\mycsreg/_0613_ ), .Z(\srccs_raw [2] ) );
BUF_X1 \mycsreg/_1585_ ( .A(\mycsreg/CSReg[3][3] ), .Z(\mycsreg/_0121_ ) );
BUF_X1 \mycsreg/_1586_ ( .A(\mycsreg/CSReg[2][3] ), .Z(\mycsreg/_0089_ ) );
BUF_X1 \mycsreg/_1587_ ( .A(\mycsreg/CSReg[1][3] ), .Z(\mycsreg/_0057_ ) );
BUF_X1 \mycsreg/_1588_ ( .A(\mycsreg/CSReg[0][3] ), .Z(\mycsreg/_0025_ ) );
BUF_X1 \mycsreg/_1589_ ( .A(\mycsreg/_0616_ ), .Z(\srccs_raw [3] ) );
BUF_X1 \mycsreg/_1590_ ( .A(\mycsreg/CSReg[3][4] ), .Z(\mycsreg/_0122_ ) );
BUF_X1 \mycsreg/_1591_ ( .A(\mycsreg/CSReg[2][4] ), .Z(\mycsreg/_0090_ ) );
BUF_X1 \mycsreg/_1592_ ( .A(\mycsreg/CSReg[1][4] ), .Z(\mycsreg/_0058_ ) );
BUF_X1 \mycsreg/_1593_ ( .A(\mycsreg/CSReg[0][4] ), .Z(\mycsreg/_0026_ ) );
BUF_X1 \mycsreg/_1594_ ( .A(\mycsreg/_0617_ ), .Z(\srccs_raw [4] ) );
BUF_X1 \mycsreg/_1595_ ( .A(\mycsreg/CSReg[3][5] ), .Z(\mycsreg/_0123_ ) );
BUF_X1 \mycsreg/_1596_ ( .A(\mycsreg/CSReg[2][5] ), .Z(\mycsreg/_0091_ ) );
BUF_X1 \mycsreg/_1597_ ( .A(\mycsreg/CSReg[1][5] ), .Z(\mycsreg/_0059_ ) );
BUF_X1 \mycsreg/_1598_ ( .A(\mycsreg/CSReg[0][5] ), .Z(\mycsreg/_0027_ ) );
BUF_X1 \mycsreg/_1599_ ( .A(\mycsreg/_0618_ ), .Z(\srccs_raw [5] ) );
BUF_X1 \mycsreg/_1600_ ( .A(\mycsreg/CSReg[3][6] ), .Z(\mycsreg/_0124_ ) );
BUF_X1 \mycsreg/_1601_ ( .A(\mycsreg/CSReg[2][6] ), .Z(\mycsreg/_0092_ ) );
BUF_X1 \mycsreg/_1602_ ( .A(\mycsreg/CSReg[1][6] ), .Z(\mycsreg/_0060_ ) );
BUF_X1 \mycsreg/_1603_ ( .A(\mycsreg/CSReg[0][6] ), .Z(\mycsreg/_0028_ ) );
BUF_X1 \mycsreg/_1604_ ( .A(\mycsreg/_0619_ ), .Z(\srccs_raw [6] ) );
BUF_X1 \mycsreg/_1605_ ( .A(\mycsreg/CSReg[3][7] ), .Z(\mycsreg/_0125_ ) );
BUF_X1 \mycsreg/_1606_ ( .A(\mycsreg/CSReg[2][7] ), .Z(\mycsreg/_0093_ ) );
BUF_X1 \mycsreg/_1607_ ( .A(\mycsreg/CSReg[1][7] ), .Z(\mycsreg/_0061_ ) );
BUF_X1 \mycsreg/_1608_ ( .A(\mycsreg/CSReg[0][7] ), .Z(\mycsreg/_0029_ ) );
BUF_X1 \mycsreg/_1609_ ( .A(\mycsreg/_0620_ ), .Z(\srccs_raw [7] ) );
BUF_X1 \mycsreg/_1610_ ( .A(\mycsreg/CSReg[3][8] ), .Z(\mycsreg/_0126_ ) );
BUF_X1 \mycsreg/_1611_ ( .A(\mycsreg/CSReg[2][8] ), .Z(\mycsreg/_0094_ ) );
BUF_X1 \mycsreg/_1612_ ( .A(\mycsreg/CSReg[1][8] ), .Z(\mycsreg/_0062_ ) );
BUF_X1 \mycsreg/_1613_ ( .A(\mycsreg/CSReg[0][8] ), .Z(\mycsreg/_0030_ ) );
BUF_X1 \mycsreg/_1614_ ( .A(\mycsreg/_0621_ ), .Z(\srccs_raw [8] ) );
BUF_X1 \mycsreg/_1615_ ( .A(\mycsreg/CSReg[3][9] ), .Z(\mycsreg/_0127_ ) );
BUF_X1 \mycsreg/_1616_ ( .A(\mycsreg/CSReg[2][9] ), .Z(\mycsreg/_0095_ ) );
BUF_X1 \mycsreg/_1617_ ( .A(\mycsreg/CSReg[1][9] ), .Z(\mycsreg/_0063_ ) );
BUF_X1 \mycsreg/_1618_ ( .A(\mycsreg/CSReg[0][9] ), .Z(\mycsreg/_0031_ ) );
BUF_X1 \mycsreg/_1619_ ( .A(\mycsreg/_0622_ ), .Z(\srccs_raw [9] ) );
BUF_X1 \mycsreg/_1620_ ( .A(\mycsreg/CSReg[3][10] ), .Z(\mycsreg/_0097_ ) );
BUF_X1 \mycsreg/_1621_ ( .A(\mycsreg/CSReg[2][10] ), .Z(\mycsreg/_0065_ ) );
BUF_X1 \mycsreg/_1622_ ( .A(\mycsreg/CSReg[1][10] ), .Z(\mycsreg/_0033_ ) );
BUF_X1 \mycsreg/_1623_ ( .A(\mycsreg/CSReg[0][10] ), .Z(\mycsreg/_0001_ ) );
BUF_X1 \mycsreg/_1624_ ( .A(\mycsreg/_0592_ ), .Z(\srccs_raw [10] ) );
BUF_X1 \mycsreg/_1625_ ( .A(\mycsreg/CSReg[3][11] ), .Z(\mycsreg/_0098_ ) );
BUF_X1 \mycsreg/_1626_ ( .A(\mycsreg/CSReg[2][11] ), .Z(\mycsreg/_0066_ ) );
BUF_X1 \mycsreg/_1627_ ( .A(\mycsreg/CSReg[1][11] ), .Z(\mycsreg/_0034_ ) );
BUF_X1 \mycsreg/_1628_ ( .A(\mycsreg/CSReg[0][11] ), .Z(\mycsreg/_0002_ ) );
BUF_X1 \mycsreg/_1629_ ( .A(\mycsreg/_0593_ ), .Z(\srccs_raw [11] ) );
BUF_X1 \mycsreg/_1630_ ( .A(\mycsreg/CSReg[3][12] ), .Z(\mycsreg/_0099_ ) );
BUF_X1 \mycsreg/_1631_ ( .A(\mycsreg/CSReg[2][12] ), .Z(\mycsreg/_0067_ ) );
BUF_X1 \mycsreg/_1632_ ( .A(\mycsreg/CSReg[1][12] ), .Z(\mycsreg/_0035_ ) );
BUF_X1 \mycsreg/_1633_ ( .A(\mycsreg/CSReg[0][12] ), .Z(\mycsreg/_0003_ ) );
BUF_X1 \mycsreg/_1634_ ( .A(\mycsreg/_0594_ ), .Z(\srccs_raw [12] ) );
BUF_X1 \mycsreg/_1635_ ( .A(\mycsreg/CSReg[3][13] ), .Z(\mycsreg/_0100_ ) );
BUF_X1 \mycsreg/_1636_ ( .A(\mycsreg/CSReg[2][13] ), .Z(\mycsreg/_0068_ ) );
BUF_X1 \mycsreg/_1637_ ( .A(\mycsreg/CSReg[1][13] ), .Z(\mycsreg/_0036_ ) );
BUF_X1 \mycsreg/_1638_ ( .A(\mycsreg/CSReg[0][13] ), .Z(\mycsreg/_0004_ ) );
BUF_X1 \mycsreg/_1639_ ( .A(\mycsreg/_0595_ ), .Z(\srccs_raw [13] ) );
BUF_X1 \mycsreg/_1640_ ( .A(\mycsreg/CSReg[3][14] ), .Z(\mycsreg/_0101_ ) );
BUF_X1 \mycsreg/_1641_ ( .A(\mycsreg/CSReg[2][14] ), .Z(\mycsreg/_0069_ ) );
BUF_X1 \mycsreg/_1642_ ( .A(\mycsreg/CSReg[1][14] ), .Z(\mycsreg/_0037_ ) );
BUF_X1 \mycsreg/_1643_ ( .A(\mycsreg/CSReg[0][14] ), .Z(\mycsreg/_0005_ ) );
BUF_X1 \mycsreg/_1644_ ( .A(\mycsreg/_0596_ ), .Z(\srccs_raw [14] ) );
BUF_X1 \mycsreg/_1645_ ( .A(\mycsreg/CSReg[3][15] ), .Z(\mycsreg/_0102_ ) );
BUF_X1 \mycsreg/_1646_ ( .A(\mycsreg/CSReg[2][15] ), .Z(\mycsreg/_0070_ ) );
BUF_X1 \mycsreg/_1647_ ( .A(\mycsreg/CSReg[1][15] ), .Z(\mycsreg/_0038_ ) );
BUF_X1 \mycsreg/_1648_ ( .A(\mycsreg/CSReg[0][15] ), .Z(\mycsreg/_0006_ ) );
BUF_X1 \mycsreg/_1649_ ( .A(\mycsreg/_0597_ ), .Z(\srccs_raw [15] ) );
BUF_X1 \mycsreg/_1650_ ( .A(\mycsreg/CSReg[3][16] ), .Z(\mycsreg/_0103_ ) );
BUF_X1 \mycsreg/_1651_ ( .A(\mycsreg/CSReg[2][16] ), .Z(\mycsreg/_0071_ ) );
BUF_X1 \mycsreg/_1652_ ( .A(\mycsreg/CSReg[1][16] ), .Z(\mycsreg/_0039_ ) );
BUF_X1 \mycsreg/_1653_ ( .A(\mycsreg/CSReg[0][16] ), .Z(\mycsreg/_0007_ ) );
BUF_X1 \mycsreg/_1654_ ( .A(\mycsreg/_0598_ ), .Z(\srccs_raw [16] ) );
BUF_X1 \mycsreg/_1655_ ( .A(\mycsreg/CSReg[3][17] ), .Z(\mycsreg/_0104_ ) );
BUF_X1 \mycsreg/_1656_ ( .A(\mycsreg/CSReg[2][17] ), .Z(\mycsreg/_0072_ ) );
BUF_X1 \mycsreg/_1657_ ( .A(\mycsreg/CSReg[1][17] ), .Z(\mycsreg/_0040_ ) );
BUF_X1 \mycsreg/_1658_ ( .A(\mycsreg/CSReg[0][17] ), .Z(\mycsreg/_0008_ ) );
BUF_X1 \mycsreg/_1659_ ( .A(\mycsreg/_0599_ ), .Z(\srccs_raw [17] ) );
BUF_X1 \mycsreg/_1660_ ( .A(\mycsreg/CSReg[3][18] ), .Z(\mycsreg/_0105_ ) );
BUF_X1 \mycsreg/_1661_ ( .A(\mycsreg/CSReg[2][18] ), .Z(\mycsreg/_0073_ ) );
BUF_X1 \mycsreg/_1662_ ( .A(\mycsreg/CSReg[1][18] ), .Z(\mycsreg/_0041_ ) );
BUF_X1 \mycsreg/_1663_ ( .A(\mycsreg/CSReg[0][18] ), .Z(\mycsreg/_0009_ ) );
BUF_X1 \mycsreg/_1664_ ( .A(\mycsreg/_0600_ ), .Z(\srccs_raw [18] ) );
BUF_X1 \mycsreg/_1665_ ( .A(\mycsreg/CSReg[3][19] ), .Z(\mycsreg/_0106_ ) );
BUF_X1 \mycsreg/_1666_ ( .A(\mycsreg/CSReg[2][19] ), .Z(\mycsreg/_0074_ ) );
BUF_X1 \mycsreg/_1667_ ( .A(\mycsreg/CSReg[1][19] ), .Z(\mycsreg/_0042_ ) );
BUF_X1 \mycsreg/_1668_ ( .A(\mycsreg/CSReg[0][19] ), .Z(\mycsreg/_0010_ ) );
BUF_X1 \mycsreg/_1669_ ( .A(\mycsreg/_0601_ ), .Z(\srccs_raw [19] ) );
BUF_X1 \mycsreg/_1670_ ( .A(\mycsreg/CSReg[3][20] ), .Z(\mycsreg/_0108_ ) );
BUF_X1 \mycsreg/_1671_ ( .A(\mycsreg/CSReg[2][20] ), .Z(\mycsreg/_0076_ ) );
BUF_X1 \mycsreg/_1672_ ( .A(\mycsreg/CSReg[1][20] ), .Z(\mycsreg/_0044_ ) );
BUF_X1 \mycsreg/_1673_ ( .A(\mycsreg/CSReg[0][20] ), .Z(\mycsreg/_0012_ ) );
BUF_X1 \mycsreg/_1674_ ( .A(\mycsreg/_0603_ ), .Z(\srccs_raw [20] ) );
BUF_X1 \mycsreg/_1675_ ( .A(\mycsreg/CSReg[3][21] ), .Z(\mycsreg/_0109_ ) );
BUF_X1 \mycsreg/_1676_ ( .A(\mycsreg/CSReg[2][21] ), .Z(\mycsreg/_0077_ ) );
BUF_X1 \mycsreg/_1677_ ( .A(\mycsreg/CSReg[1][21] ), .Z(\mycsreg/_0045_ ) );
BUF_X1 \mycsreg/_1678_ ( .A(\mycsreg/CSReg[0][21] ), .Z(\mycsreg/_0013_ ) );
BUF_X1 \mycsreg/_1679_ ( .A(\mycsreg/_0604_ ), .Z(\srccs_raw [21] ) );
BUF_X1 \mycsreg/_1680_ ( .A(\mycsreg/CSReg[3][22] ), .Z(\mycsreg/_0110_ ) );
BUF_X1 \mycsreg/_1681_ ( .A(\mycsreg/CSReg[2][22] ), .Z(\mycsreg/_0078_ ) );
BUF_X1 \mycsreg/_1682_ ( .A(\mycsreg/CSReg[1][22] ), .Z(\mycsreg/_0046_ ) );
BUF_X1 \mycsreg/_1683_ ( .A(\mycsreg/CSReg[0][22] ), .Z(\mycsreg/_0014_ ) );
BUF_X1 \mycsreg/_1684_ ( .A(\mycsreg/_0605_ ), .Z(\srccs_raw [22] ) );
BUF_X1 \mycsreg/_1685_ ( .A(\mycsreg/CSReg[3][23] ), .Z(\mycsreg/_0111_ ) );
BUF_X1 \mycsreg/_1686_ ( .A(\mycsreg/CSReg[2][23] ), .Z(\mycsreg/_0079_ ) );
BUF_X1 \mycsreg/_1687_ ( .A(\mycsreg/CSReg[1][23] ), .Z(\mycsreg/_0047_ ) );
BUF_X1 \mycsreg/_1688_ ( .A(\mycsreg/CSReg[0][23] ), .Z(\mycsreg/_0015_ ) );
BUF_X1 \mycsreg/_1689_ ( .A(\mycsreg/_0606_ ), .Z(\srccs_raw [23] ) );
BUF_X1 \mycsreg/_1690_ ( .A(\mycsreg/CSReg[3][24] ), .Z(\mycsreg/_0112_ ) );
BUF_X1 \mycsreg/_1691_ ( .A(\mycsreg/CSReg[2][24] ), .Z(\mycsreg/_0080_ ) );
BUF_X1 \mycsreg/_1692_ ( .A(\mycsreg/CSReg[1][24] ), .Z(\mycsreg/_0048_ ) );
BUF_X1 \mycsreg/_1693_ ( .A(\mycsreg/CSReg[0][24] ), .Z(\mycsreg/_0016_ ) );
BUF_X1 \mycsreg/_1694_ ( .A(\mycsreg/_0607_ ), .Z(\srccs_raw [24] ) );
BUF_X1 \mycsreg/_1695_ ( .A(\mycsreg/CSReg[3][25] ), .Z(\mycsreg/_0113_ ) );
BUF_X1 \mycsreg/_1696_ ( .A(\mycsreg/CSReg[2][25] ), .Z(\mycsreg/_0081_ ) );
BUF_X1 \mycsreg/_1697_ ( .A(\mycsreg/CSReg[1][25] ), .Z(\mycsreg/_0049_ ) );
BUF_X1 \mycsreg/_1698_ ( .A(\mycsreg/CSReg[0][25] ), .Z(\mycsreg/_0017_ ) );
BUF_X1 \mycsreg/_1699_ ( .A(\mycsreg/_0608_ ), .Z(\srccs_raw [25] ) );
BUF_X1 \mycsreg/_1700_ ( .A(\mycsreg/CSReg[3][26] ), .Z(\mycsreg/_0114_ ) );
BUF_X1 \mycsreg/_1701_ ( .A(\mycsreg/CSReg[2][26] ), .Z(\mycsreg/_0082_ ) );
BUF_X1 \mycsreg/_1702_ ( .A(\mycsreg/CSReg[1][26] ), .Z(\mycsreg/_0050_ ) );
BUF_X1 \mycsreg/_1703_ ( .A(\mycsreg/CSReg[0][26] ), .Z(\mycsreg/_0018_ ) );
BUF_X1 \mycsreg/_1704_ ( .A(\mycsreg/_0609_ ), .Z(\srccs_raw [26] ) );
BUF_X1 \mycsreg/_1705_ ( .A(\mycsreg/CSReg[3][27] ), .Z(\mycsreg/_0115_ ) );
BUF_X1 \mycsreg/_1706_ ( .A(\mycsreg/CSReg[2][27] ), .Z(\mycsreg/_0083_ ) );
BUF_X1 \mycsreg/_1707_ ( .A(\mycsreg/CSReg[1][27] ), .Z(\mycsreg/_0051_ ) );
BUF_X1 \mycsreg/_1708_ ( .A(\mycsreg/CSReg[0][27] ), .Z(\mycsreg/_0019_ ) );
BUF_X1 \mycsreg/_1709_ ( .A(\mycsreg/_0610_ ), .Z(\srccs_raw [27] ) );
BUF_X1 \mycsreg/_1710_ ( .A(\mycsreg/CSReg[3][28] ), .Z(\mycsreg/_0116_ ) );
BUF_X1 \mycsreg/_1711_ ( .A(\mycsreg/CSReg[2][28] ), .Z(\mycsreg/_0084_ ) );
BUF_X1 \mycsreg/_1712_ ( .A(\mycsreg/CSReg[1][28] ), .Z(\mycsreg/_0052_ ) );
BUF_X1 \mycsreg/_1713_ ( .A(\mycsreg/CSReg[0][28] ), .Z(\mycsreg/_0020_ ) );
BUF_X1 \mycsreg/_1714_ ( .A(\mycsreg/_0611_ ), .Z(\srccs_raw [28] ) );
BUF_X1 \mycsreg/_1715_ ( .A(\mycsreg/CSReg[3][29] ), .Z(\mycsreg/_0117_ ) );
BUF_X1 \mycsreg/_1716_ ( .A(\mycsreg/CSReg[2][29] ), .Z(\mycsreg/_0085_ ) );
BUF_X1 \mycsreg/_1717_ ( .A(\mycsreg/CSReg[1][29] ), .Z(\mycsreg/_0053_ ) );
BUF_X1 \mycsreg/_1718_ ( .A(\mycsreg/CSReg[0][29] ), .Z(\mycsreg/_0021_ ) );
BUF_X1 \mycsreg/_1719_ ( .A(\mycsreg/_0612_ ), .Z(\srccs_raw [29] ) );
BUF_X1 \mycsreg/_1720_ ( .A(\mycsreg/CSReg[3][30] ), .Z(\mycsreg/_0119_ ) );
BUF_X1 \mycsreg/_1721_ ( .A(\mycsreg/CSReg[2][30] ), .Z(\mycsreg/_0087_ ) );
BUF_X1 \mycsreg/_1722_ ( .A(\mycsreg/CSReg[1][30] ), .Z(\mycsreg/_0055_ ) );
BUF_X1 \mycsreg/_1723_ ( .A(\mycsreg/CSReg[0][30] ), .Z(\mycsreg/_0023_ ) );
BUF_X1 \mycsreg/_1724_ ( .A(\mycsreg/_0614_ ), .Z(\srccs_raw [30] ) );
BUF_X1 \mycsreg/_1725_ ( .A(\mycsreg/CSReg[3][31] ), .Z(\mycsreg/_0120_ ) );
BUF_X1 \mycsreg/_1726_ ( .A(\mycsreg/CSReg[2][31] ), .Z(\mycsreg/_0088_ ) );
BUF_X1 \mycsreg/_1727_ ( .A(\mycsreg/CSReg[1][31] ), .Z(\mycsreg/_0056_ ) );
BUF_X1 \mycsreg/_1728_ ( .A(\mycsreg/CSReg[0][31] ), .Z(\mycsreg/_0024_ ) );
BUF_X1 \mycsreg/_1729_ ( .A(\mycsreg/_0615_ ), .Z(\srccs_raw [31] ) );
BUF_X1 \mycsreg/_1730_ ( .A(\LS_WB_wdata_csreg [0] ), .Z(\mycsreg/_0636_ ) );
BUF_X1 \mycsreg/_1731_ ( .A(\LS_WB_wen_csreg [0] ), .Z(\mycsreg/_0668_ ) );
BUF_X1 \mycsreg/_1732_ ( .A(\LS_WB_wdata_csreg [1] ), .Z(\mycsreg/_0647_ ) );
BUF_X1 \mycsreg/_1733_ ( .A(\LS_WB_wen_csreg [1] ), .Z(\mycsreg/_0669_ ) );
BUF_X1 \mycsreg/_1734_ ( .A(\LS_WB_wdata_csreg [2] ), .Z(\mycsreg/_0658_ ) );
BUF_X1 \mycsreg/_1735_ ( .A(\LS_WB_wen_csreg [2] ), .Z(\mycsreg/_0670_ ) );
BUF_X1 \mycsreg/_1736_ ( .A(\LS_WB_wdata_csreg [3] ), .Z(\mycsreg/_0661_ ) );
BUF_X1 \mycsreg/_1737_ ( .A(\LS_WB_wen_csreg [3] ), .Z(\mycsreg/_0671_ ) );
BUF_X1 \mycsreg/_1738_ ( .A(\LS_WB_wdata_csreg [4] ), .Z(\mycsreg/_0662_ ) );
BUF_X1 \mycsreg/_1739_ ( .A(\LS_WB_wen_csreg [4] ), .Z(\mycsreg/_0672_ ) );
BUF_X1 \mycsreg/_1740_ ( .A(\LS_WB_wdata_csreg [5] ), .Z(\mycsreg/_0663_ ) );
BUF_X1 \mycsreg/_1741_ ( .A(\LS_WB_wen_csreg [5] ), .Z(\mycsreg/_0673_ ) );
BUF_X1 \mycsreg/_1742_ ( .A(\mycsreg/_0128_ ), .Z(\mycsreg/_0804_ ) );
BUF_X1 \mycsreg/_1743_ ( .A(\mycsreg/_0129_ ), .Z(\mycsreg/_0805_ ) );
BUF_X1 \mycsreg/_1744_ ( .A(\mycsreg/_0130_ ), .Z(\mycsreg/_0806_ ) );
BUF_X1 \mycsreg/_1745_ ( .A(\mycsreg/_0131_ ), .Z(\mycsreg/_0807_ ) );
BUF_X1 \mycsreg/_1746_ ( .A(\mycsreg/_0132_ ), .Z(\mycsreg/_0808_ ) );
BUF_X1 \mycsreg/_1747_ ( .A(\mycsreg/_0133_ ), .Z(\mycsreg/_0809_ ) );
BUF_X1 \mycsreg/_1748_ ( .A(\mycsreg/_0134_ ), .Z(\mycsreg/_0810_ ) );
BUF_X1 \mycsreg/_1749_ ( .A(\mycsreg/_0135_ ), .Z(\mycsreg/_0811_ ) );
BUF_X1 \mycsreg/_1750_ ( .A(\mycsreg/_0136_ ), .Z(\mycsreg/_0812_ ) );
BUF_X1 \mycsreg/_1751_ ( .A(\mycsreg/_0137_ ), .Z(\mycsreg/_0813_ ) );
BUF_X1 \mycsreg/_1752_ ( .A(\mycsreg/_0138_ ), .Z(\mycsreg/_0814_ ) );
BUF_X1 \mycsreg/_1753_ ( .A(\mycsreg/_0139_ ), .Z(\mycsreg/_0815_ ) );
BUF_X1 \mycsreg/_1754_ ( .A(\LS_WB_wdata_csreg [6] ), .Z(\mycsreg/_0664_ ) );
BUF_X1 \mycsreg/_1755_ ( .A(\mycsreg/_0140_ ), .Z(\mycsreg/_0816_ ) );
BUF_X1 \mycsreg/_1756_ ( .A(\LS_WB_wdata_csreg [7] ), .Z(\mycsreg/_0665_ ) );
BUF_X1 \mycsreg/_1757_ ( .A(\mycsreg/_0141_ ), .Z(\mycsreg/_0817_ ) );
BUF_X1 \mycsreg/_1758_ ( .A(\LS_WB_wdata_csreg [8] ), .Z(\mycsreg/_0666_ ) );
BUF_X1 \mycsreg/_1759_ ( .A(\mycsreg/_0142_ ), .Z(\mycsreg/_0818_ ) );
BUF_X1 \mycsreg/_1760_ ( .A(\LS_WB_wdata_csreg [9] ), .Z(\mycsreg/_0667_ ) );
BUF_X1 \mycsreg/_1761_ ( .A(\mycsreg/_0143_ ), .Z(\mycsreg/_0819_ ) );
BUF_X1 \mycsreg/_1762_ ( .A(\LS_WB_wdata_csreg [10] ), .Z(\mycsreg/_0637_ ) );
BUF_X1 \mycsreg/_1763_ ( .A(\mycsreg/_0144_ ), .Z(\mycsreg/_0820_ ) );
BUF_X1 \mycsreg/_1764_ ( .A(\LS_WB_wdata_csreg [11] ), .Z(\mycsreg/_0638_ ) );
BUF_X1 \mycsreg/_1765_ ( .A(\mycsreg/_0145_ ), .Z(\mycsreg/_0821_ ) );
BUF_X1 \mycsreg/_1766_ ( .A(\LS_WB_wdata_csreg [12] ), .Z(\mycsreg/_0639_ ) );
BUF_X1 \mycsreg/_1767_ ( .A(\mycsreg/_0146_ ), .Z(\mycsreg/_0822_ ) );
BUF_X1 \mycsreg/_1768_ ( .A(\LS_WB_wdata_csreg [13] ), .Z(\mycsreg/_0640_ ) );
BUF_X1 \mycsreg/_1769_ ( .A(\mycsreg/_0147_ ), .Z(\mycsreg/_0823_ ) );
BUF_X1 \mycsreg/_1770_ ( .A(\LS_WB_wdata_csreg [14] ), .Z(\mycsreg/_0641_ ) );
BUF_X1 \mycsreg/_1771_ ( .A(\mycsreg/_0148_ ), .Z(\mycsreg/_0824_ ) );
BUF_X1 \mycsreg/_1772_ ( .A(\LS_WB_wdata_csreg [15] ), .Z(\mycsreg/_0642_ ) );
BUF_X1 \mycsreg/_1773_ ( .A(\mycsreg/_0149_ ), .Z(\mycsreg/_0825_ ) );
BUF_X1 \mycsreg/_1774_ ( .A(\LS_WB_wdata_csreg [16] ), .Z(\mycsreg/_0643_ ) );
BUF_X1 \mycsreg/_1775_ ( .A(\mycsreg/_0150_ ), .Z(\mycsreg/_0826_ ) );
BUF_X1 \mycsreg/_1776_ ( .A(\LS_WB_wdata_csreg [17] ), .Z(\mycsreg/_0644_ ) );
BUF_X1 \mycsreg/_1777_ ( .A(\mycsreg/_0151_ ), .Z(\mycsreg/_0827_ ) );
BUF_X1 \mycsreg/_1778_ ( .A(\LS_WB_wdata_csreg [18] ), .Z(\mycsreg/_0645_ ) );
BUF_X1 \mycsreg/_1779_ ( .A(\mycsreg/_0152_ ), .Z(\mycsreg/_0828_ ) );
BUF_X1 \mycsreg/_1780_ ( .A(\LS_WB_wdata_csreg [19] ), .Z(\mycsreg/_0646_ ) );
BUF_X1 \mycsreg/_1781_ ( .A(\mycsreg/_0153_ ), .Z(\mycsreg/_0829_ ) );
BUF_X1 \mycsreg/_1782_ ( .A(\LS_WB_wdata_csreg [20] ), .Z(\mycsreg/_0648_ ) );
BUF_X1 \mycsreg/_1783_ ( .A(\mycsreg/_0154_ ), .Z(\mycsreg/_0830_ ) );
BUF_X1 \mycsreg/_1784_ ( .A(\LS_WB_wdata_csreg [21] ), .Z(\mycsreg/_0649_ ) );
BUF_X1 \mycsreg/_1785_ ( .A(\mycsreg/_0155_ ), .Z(\mycsreg/_0831_ ) );
BUF_X1 \mycsreg/_1786_ ( .A(\LS_WB_wdata_csreg [22] ), .Z(\mycsreg/_0650_ ) );
BUF_X1 \mycsreg/_1787_ ( .A(\mycsreg/_0156_ ), .Z(\mycsreg/_0832_ ) );
BUF_X1 \mycsreg/_1788_ ( .A(\LS_WB_wdata_csreg [23] ), .Z(\mycsreg/_0651_ ) );
BUF_X1 \mycsreg/_1789_ ( .A(\mycsreg/_0157_ ), .Z(\mycsreg/_0833_ ) );
BUF_X1 \mycsreg/_1790_ ( .A(\LS_WB_wdata_csreg [24] ), .Z(\mycsreg/_0652_ ) );
BUF_X1 \mycsreg/_1791_ ( .A(\mycsreg/_0158_ ), .Z(\mycsreg/_0834_ ) );
BUF_X1 \mycsreg/_1792_ ( .A(\LS_WB_wdata_csreg [25] ), .Z(\mycsreg/_0653_ ) );
BUF_X1 \mycsreg/_1793_ ( .A(\mycsreg/_0159_ ), .Z(\mycsreg/_0835_ ) );
BUF_X1 \mycsreg/_1794_ ( .A(\LS_WB_wdata_csreg [26] ), .Z(\mycsreg/_0654_ ) );
BUF_X1 \mycsreg/_1795_ ( .A(\mycsreg/_0160_ ), .Z(\mycsreg/_0836_ ) );
BUF_X1 \mycsreg/_1796_ ( .A(\LS_WB_wdata_csreg [27] ), .Z(\mycsreg/_0655_ ) );
BUF_X1 \mycsreg/_1797_ ( .A(\mycsreg/_0161_ ), .Z(\mycsreg/_0837_ ) );
BUF_X1 \mycsreg/_1798_ ( .A(\LS_WB_wdata_csreg [28] ), .Z(\mycsreg/_0656_ ) );
BUF_X1 \mycsreg/_1799_ ( .A(\mycsreg/_0162_ ), .Z(\mycsreg/_0838_ ) );
BUF_X1 \mycsreg/_1800_ ( .A(\LS_WB_wdata_csreg [29] ), .Z(\mycsreg/_0657_ ) );
BUF_X1 \mycsreg/_1801_ ( .A(\mycsreg/_0163_ ), .Z(\mycsreg/_0839_ ) );
BUF_X1 \mycsreg/_1802_ ( .A(\LS_WB_wdata_csreg [30] ), .Z(\mycsreg/_0659_ ) );
BUF_X1 \mycsreg/_1803_ ( .A(\mycsreg/_0164_ ), .Z(\mycsreg/_0840_ ) );
BUF_X1 \mycsreg/_1804_ ( .A(\LS_WB_wdata_csreg [31] ), .Z(\mycsreg/_0660_ ) );
BUF_X1 \mycsreg/_1805_ ( .A(\mycsreg/_0165_ ), .Z(\mycsreg/_0841_ ) );
BUF_X1 \mycsreg/_1806_ ( .A(\mycsreg/_0166_ ), .Z(\mycsreg/_0842_ ) );
BUF_X1 \mycsreg/_1807_ ( .A(\mycsreg/_0167_ ), .Z(\mycsreg/_0843_ ) );
BUF_X1 \mycsreg/_1808_ ( .A(\mycsreg/_0168_ ), .Z(\mycsreg/_0844_ ) );
BUF_X1 \mycsreg/_1809_ ( .A(\mycsreg/_0169_ ), .Z(\mycsreg/_0845_ ) );
BUF_X1 \mycsreg/_1810_ ( .A(\mycsreg/_0170_ ), .Z(\mycsreg/_0846_ ) );
BUF_X1 \mycsreg/_1811_ ( .A(\mycsreg/_0171_ ), .Z(\mycsreg/_0847_ ) );
BUF_X1 \mycsreg/_1812_ ( .A(\mycsreg/_0172_ ), .Z(\mycsreg/_0848_ ) );
BUF_X1 \mycsreg/_1813_ ( .A(\mycsreg/_0173_ ), .Z(\mycsreg/_0849_ ) );
BUF_X1 \mycsreg/_1814_ ( .A(\mycsreg/_0174_ ), .Z(\mycsreg/_0850_ ) );
BUF_X1 \mycsreg/_1815_ ( .A(\mycsreg/_0175_ ), .Z(\mycsreg/_0851_ ) );
BUF_X1 \mycsreg/_1816_ ( .A(\mycsreg/_0176_ ), .Z(\mycsreg/_0852_ ) );
BUF_X1 \mycsreg/_1817_ ( .A(\mycsreg/_0177_ ), .Z(\mycsreg/_0853_ ) );
BUF_X1 \mycsreg/_1818_ ( .A(\mycsreg/_0178_ ), .Z(\mycsreg/_0854_ ) );
BUF_X1 \mycsreg/_1819_ ( .A(\mycsreg/_0179_ ), .Z(\mycsreg/_0855_ ) );
BUF_X1 \mycsreg/_1820_ ( .A(\mycsreg/_0180_ ), .Z(\mycsreg/_0856_ ) );
BUF_X1 \mycsreg/_1821_ ( .A(\mycsreg/_0181_ ), .Z(\mycsreg/_0857_ ) );
BUF_X1 \mycsreg/_1822_ ( .A(\mycsreg/_0182_ ), .Z(\mycsreg/_0858_ ) );
BUF_X1 \mycsreg/_1823_ ( .A(\mycsreg/_0183_ ), .Z(\mycsreg/_0859_ ) );
BUF_X1 \mycsreg/_1824_ ( .A(\mycsreg/_0184_ ), .Z(\mycsreg/_0860_ ) );
BUF_X1 \mycsreg/_1825_ ( .A(\mycsreg/_0185_ ), .Z(\mycsreg/_0861_ ) );
BUF_X1 \mycsreg/_1826_ ( .A(\mycsreg/_0186_ ), .Z(\mycsreg/_0862_ ) );
BUF_X1 \mycsreg/_1827_ ( .A(\mycsreg/_0187_ ), .Z(\mycsreg/_0863_ ) );
BUF_X1 \mycsreg/_1828_ ( .A(\mycsreg/_0188_ ), .Z(\mycsreg/_0864_ ) );
BUF_X1 \mycsreg/_1829_ ( .A(\mycsreg/_0189_ ), .Z(\mycsreg/_0865_ ) );
BUF_X1 \mycsreg/_1830_ ( .A(\mycsreg/_0190_ ), .Z(\mycsreg/_0866_ ) );
BUF_X1 \mycsreg/_1831_ ( .A(\mycsreg/_0191_ ), .Z(\mycsreg/_0867_ ) );
BUF_X1 \mycsreg/_1832_ ( .A(\mycsreg/_0192_ ), .Z(\mycsreg/_0868_ ) );
BUF_X1 \mycsreg/_1833_ ( .A(\mycsreg/_0193_ ), .Z(\mycsreg/_0869_ ) );
BUF_X1 \mycsreg/_1834_ ( .A(\mycsreg/_0194_ ), .Z(\mycsreg/_0870_ ) );
BUF_X1 \mycsreg/_1835_ ( .A(\mycsreg/_0195_ ), .Z(\mycsreg/_0871_ ) );
BUF_X1 \mycsreg/_1836_ ( .A(\mycsreg/_0196_ ), .Z(\mycsreg/_0872_ ) );
BUF_X1 \mycsreg/_1837_ ( .A(\mycsreg/_0197_ ), .Z(\mycsreg/_0873_ ) );
BUF_X1 \mycsreg/_1838_ ( .A(\mycsreg/_0198_ ), .Z(\mycsreg/_0874_ ) );
BUF_X1 \mycsreg/_1839_ ( .A(\mycsreg/_0199_ ), .Z(\mycsreg/_0875_ ) );
BUF_X1 \mycsreg/_1840_ ( .A(\mycsreg/_0200_ ), .Z(\mycsreg/_0876_ ) );
BUF_X1 \mycsreg/_1841_ ( .A(\mycsreg/_0201_ ), .Z(\mycsreg/_0877_ ) );
BUF_X1 \mycsreg/_1842_ ( .A(\mycsreg/_0202_ ), .Z(\mycsreg/_0878_ ) );
BUF_X1 \mycsreg/_1843_ ( .A(\mycsreg/_0203_ ), .Z(\mycsreg/_0879_ ) );
BUF_X1 \mycsreg/_1844_ ( .A(\mycsreg/_0204_ ), .Z(\mycsreg/_0880_ ) );
BUF_X1 \mycsreg/_1845_ ( .A(\mycsreg/_0205_ ), .Z(\mycsreg/_0881_ ) );
BUF_X1 \mycsreg/_1846_ ( .A(\mycsreg/_0206_ ), .Z(\mycsreg/_0882_ ) );
BUF_X1 \mycsreg/_1847_ ( .A(\mycsreg/_0207_ ), .Z(\mycsreg/_0883_ ) );
BUF_X1 \mycsreg/_1848_ ( .A(\mycsreg/_0208_ ), .Z(\mycsreg/_0884_ ) );
BUF_X1 \mycsreg/_1849_ ( .A(\mycsreg/_0209_ ), .Z(\mycsreg/_0885_ ) );
BUF_X1 \mycsreg/_1850_ ( .A(\mycsreg/_0210_ ), .Z(\mycsreg/_0886_ ) );
BUF_X1 \mycsreg/_1851_ ( .A(\mycsreg/_0211_ ), .Z(\mycsreg/_0887_ ) );
BUF_X1 \mycsreg/_1852_ ( .A(\mycsreg/_0212_ ), .Z(\mycsreg/_0888_ ) );
BUF_X1 \mycsreg/_1853_ ( .A(\mycsreg/_0213_ ), .Z(\mycsreg/_0889_ ) );
BUF_X1 \mycsreg/_1854_ ( .A(\mycsreg/_0214_ ), .Z(\mycsreg/_0890_ ) );
BUF_X1 \mycsreg/_1855_ ( .A(\mycsreg/_0215_ ), .Z(\mycsreg/_0891_ ) );
BUF_X1 \mycsreg/_1856_ ( .A(\mycsreg/_0216_ ), .Z(\mycsreg/_0892_ ) );
BUF_X1 \mycsreg/_1857_ ( .A(\mycsreg/_0217_ ), .Z(\mycsreg/_0893_ ) );
BUF_X1 \mycsreg/_1858_ ( .A(\mycsreg/_0218_ ), .Z(\mycsreg/_0894_ ) );
BUF_X1 \mycsreg/_1859_ ( .A(\mycsreg/_0219_ ), .Z(\mycsreg/_0895_ ) );
BUF_X1 \mycsreg/_1860_ ( .A(\mycsreg/_0220_ ), .Z(\mycsreg/_0896_ ) );
BUF_X1 \mycsreg/_1861_ ( .A(\mycsreg/_0221_ ), .Z(\mycsreg/_0897_ ) );
BUF_X1 \mycsreg/_1862_ ( .A(\mycsreg/_0222_ ), .Z(\mycsreg/_0898_ ) );
BUF_X1 \mycsreg/_1863_ ( .A(\mycsreg/_0223_ ), .Z(\mycsreg/_0899_ ) );
BUF_X1 \mycsreg/_1864_ ( .A(\mycsreg/_0224_ ), .Z(\mycsreg/_0900_ ) );
BUF_X1 \mycsreg/_1865_ ( .A(\mycsreg/_0225_ ), .Z(\mycsreg/_0901_ ) );
BUF_X1 \mycsreg/_1866_ ( .A(\mycsreg/_0226_ ), .Z(\mycsreg/_0902_ ) );
BUF_X1 \mycsreg/_1867_ ( .A(\mycsreg/_0227_ ), .Z(\mycsreg/_0903_ ) );
BUF_X1 \mycsreg/_1868_ ( .A(\mycsreg/_0228_ ), .Z(\mycsreg/_0904_ ) );
BUF_X1 \mycsreg/_1869_ ( .A(\mycsreg/_0229_ ), .Z(\mycsreg/_0905_ ) );
BUF_X1 \mycsreg/_1870_ ( .A(\mycsreg/_0230_ ), .Z(\mycsreg/_0906_ ) );
BUF_X1 \mycsreg/_1871_ ( .A(\mycsreg/_0231_ ), .Z(\mycsreg/_0907_ ) );
BUF_X1 \mycsreg/_1872_ ( .A(\mycsreg/_0232_ ), .Z(\mycsreg/_0908_ ) );
BUF_X1 \mycsreg/_1873_ ( .A(\mycsreg/_0233_ ), .Z(\mycsreg/_0909_ ) );
BUF_X1 \mycsreg/_1874_ ( .A(\mycsreg/_0234_ ), .Z(\mycsreg/_0910_ ) );
BUF_X1 \mycsreg/_1875_ ( .A(\mycsreg/_0235_ ), .Z(\mycsreg/_0911_ ) );
BUF_X1 \mycsreg/_1876_ ( .A(\mycsreg/_0236_ ), .Z(\mycsreg/_0912_ ) );
BUF_X1 \mycsreg/_1877_ ( .A(\mycsreg/_0237_ ), .Z(\mycsreg/_0913_ ) );
BUF_X1 \mycsreg/_1878_ ( .A(\mycsreg/_0238_ ), .Z(\mycsreg/_0914_ ) );
BUF_X1 \mycsreg/_1879_ ( .A(\mycsreg/_0239_ ), .Z(\mycsreg/_0915_ ) );
BUF_X1 \mycsreg/_1880_ ( .A(\mycsreg/_0240_ ), .Z(\mycsreg/_0916_ ) );
BUF_X1 \mycsreg/_1881_ ( .A(\mycsreg/_0241_ ), .Z(\mycsreg/_0917_ ) );
BUF_X1 \mycsreg/_1882_ ( .A(\mycsreg/_0242_ ), .Z(\mycsreg/_0918_ ) );
BUF_X1 \mycsreg/_1883_ ( .A(\mycsreg/_0243_ ), .Z(\mycsreg/_0919_ ) );
BUF_X1 \mycsreg/_1884_ ( .A(\mycsreg/_0244_ ), .Z(\mycsreg/_0920_ ) );
BUF_X1 \mycsreg/_1885_ ( .A(\mycsreg/_0245_ ), .Z(\mycsreg/_0921_ ) );
BUF_X1 \mycsreg/_1886_ ( .A(\mycsreg/_0246_ ), .Z(\mycsreg/_0922_ ) );
BUF_X1 \mycsreg/_1887_ ( .A(\mycsreg/_0247_ ), .Z(\mycsreg/_0923_ ) );
BUF_X1 \mycsreg/_1888_ ( .A(\mycsreg/_0248_ ), .Z(\mycsreg/_0924_ ) );
BUF_X1 \mycsreg/_1889_ ( .A(\mycsreg/_0249_ ), .Z(\mycsreg/_0925_ ) );
BUF_X1 \mycsreg/_1890_ ( .A(\mycsreg/_0250_ ), .Z(\mycsreg/_0926_ ) );
BUF_X1 \mycsreg/_1891_ ( .A(\mycsreg/_0251_ ), .Z(\mycsreg/_0927_ ) );
BUF_X1 \mycsreg/_1892_ ( .A(\mycsreg/_0252_ ), .Z(\mycsreg/_0928_ ) );
BUF_X1 \mycsreg/_1893_ ( .A(\mycsreg/_0253_ ), .Z(\mycsreg/_0929_ ) );
BUF_X1 \mycsreg/_1894_ ( .A(\mycsreg/_0254_ ), .Z(\mycsreg/_0930_ ) );
BUF_X1 \mycsreg/_1895_ ( .A(\mycsreg/_0255_ ), .Z(\mycsreg/_0931_ ) );
MUX2_X1 \myexu/_2887_ ( .A(\myexu/_2483_ ), .B(\myexu/_0319_ ), .S(fanout_net_8 ), .Z(\myexu/_0026_ ) );
MUX2_X1 \myexu/_2888_ ( .A(\myexu/_2459_ ), .B(\myexu/_0295_ ), .S(fanout_net_8 ), .Z(\myexu/_0002_ ) );
INV_X4 \myexu/_2889_ ( .A(fanout_net_8 ), .ZN(\myexu/_1926_ ) );
NAND2_X1 \myexu/_2890_ ( .A1(\myexu/_1926_ ), .A2(\myexu/_2470_ ), .ZN(\myexu/_1927_ ) );
NAND2_X1 \myexu/_2891_ ( .A1(fanout_net_8 ), .A2(\myexu/_0306_ ), .ZN(\myexu/_1928_ ) );
NAND2_X1 \myexu/_2892_ ( .A1(\myexu/_1927_ ), .A2(\myexu/_1928_ ), .ZN(\myexu/_0013_ ) );
MUX2_X1 \myexu/_2893_ ( .A(\myexu/_2481_ ), .B(\myexu/_0317_ ), .S(fanout_net_8 ), .Z(\myexu/_0024_ ) );
INV_X2 \myexu/_2894_ ( .A(\myexu/_2484_ ), .ZN(\myexu/_1929_ ) );
NAND2_X1 \myexu/_2895_ ( .A1(\myexu/_1926_ ), .A2(\myexu/_1929_ ), .ZN(\myexu/_1930_ ) );
INV_X4 \myexu/_2896_ ( .A(\myexu/_0320_ ), .ZN(\myexu/_1931_ ) );
NAND2_X1 \myexu/_2897_ ( .A1(\myexu/_1931_ ), .A2(fanout_net_8 ), .ZN(\myexu/_1932_ ) );
AND2_X1 \myexu/_2898_ ( .A1(\myexu/_1930_ ), .A2(\myexu/_1932_ ), .ZN(\myexu/_0027_ ) );
MUX2_X1 \myexu/_2899_ ( .A(\myexu/_2485_ ), .B(\myexu/_0321_ ), .S(fanout_net_8 ), .Z(\myexu/_0028_ ) );
MUX2_X1 \myexu/_2900_ ( .A(\myexu/_2486_ ), .B(\myexu/_0322_ ), .S(fanout_net_8 ), .Z(\myexu/_0029_ ) );
MUX2_X1 \myexu/_2901_ ( .A(\myexu/_2487_ ), .B(\myexu/_0323_ ), .S(fanout_net_8 ), .Z(\myexu/_0030_ ) );
NAND2_X1 \myexu/_2902_ ( .A1(\myexu/_1926_ ), .A2(\myexu/_2488_ ), .ZN(\myexu/_1933_ ) );
NAND2_X1 \myexu/_2903_ ( .A1(fanout_net_8 ), .A2(\myexu/_0324_ ), .ZN(\myexu/_1934_ ) );
NAND2_X1 \myexu/_2904_ ( .A1(\myexu/_1933_ ), .A2(\myexu/_1934_ ), .ZN(\myexu/_0031_ ) );
MUX2_X1 \myexu/_2905_ ( .A(\myexu/_2489_ ), .B(\myexu/_0325_ ), .S(fanout_net_8 ), .Z(\myexu/_0032_ ) );
MUX2_X1 \myexu/_2906_ ( .A(\myexu/_2490_ ), .B(\myexu/_0326_ ), .S(fanout_net_8 ), .Z(\myexu/_0033_ ) );
MUX2_X1 \myexu/_2907_ ( .A(\myexu/_2460_ ), .B(\myexu/_0296_ ), .S(fanout_net_8 ), .Z(\myexu/_0003_ ) );
NAND2_X1 \myexu/_2908_ ( .A1(\myexu/_1926_ ), .A2(\myexu/_2461_ ), .ZN(\myexu/_1935_ ) );
NAND2_X1 \myexu/_2909_ ( .A1(fanout_net_8 ), .A2(\myexu/_0297_ ), .ZN(\myexu/_1936_ ) );
NAND2_X1 \myexu/_2910_ ( .A1(\myexu/_1935_ ), .A2(\myexu/_1936_ ), .ZN(\myexu/_0004_ ) );
MUX2_X1 \myexu/_2911_ ( .A(\myexu/_2462_ ), .B(\myexu/_0298_ ), .S(fanout_net_8 ), .Z(\myexu/_0005_ ) );
MUX2_X1 \myexu/_2912_ ( .A(\myexu/_2463_ ), .B(\myexu/_0299_ ), .S(fanout_net_8 ), .Z(\myexu/_0006_ ) );
MUX2_X1 \myexu/_2913_ ( .A(\myexu/_2464_ ), .B(\myexu/_0300_ ), .S(fanout_net_8 ), .Z(\myexu/_0007_ ) );
NAND2_X1 \myexu/_2914_ ( .A1(\myexu/_1926_ ), .A2(\myexu/_2465_ ), .ZN(\myexu/_1937_ ) );
NAND2_X1 \myexu/_2915_ ( .A1(fanout_net_8 ), .A2(\myexu/_0301_ ), .ZN(\myexu/_1938_ ) );
NAND2_X1 \myexu/_2916_ ( .A1(\myexu/_1937_ ), .A2(\myexu/_1938_ ), .ZN(\myexu/_0008_ ) );
BUF_X4 \myexu/_2917_ ( .A(\myexu/_1926_ ), .Z(\myexu/_1939_ ) );
NOR2_X1 \myexu/_2918_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_0302_ ), .ZN(\myexu/_1940_ ) );
NOR2_X1 \myexu/_2919_ ( .A1(fanout_net_8 ), .A2(\myexu/_2466_ ), .ZN(\myexu/_1941_ ) );
NOR2_X1 \myexu/_2920_ ( .A1(\myexu/_1940_ ), .A2(\myexu/_1941_ ), .ZN(\myexu/_0009_ ) );
NAND2_X1 \myexu/_2921_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_2467_ ), .ZN(\myexu/_1942_ ) );
NAND2_X1 \myexu/_2922_ ( .A1(fanout_net_8 ), .A2(\myexu/_0303_ ), .ZN(\myexu/_1943_ ) );
NAND2_X1 \myexu/_2923_ ( .A1(\myexu/_1942_ ), .A2(\myexu/_1943_ ), .ZN(\myexu/_0010_ ) );
MUX2_X1 \myexu/_2924_ ( .A(\myexu/_2468_ ), .B(\myexu/_0304_ ), .S(fanout_net_8 ), .Z(\myexu/_0011_ ) );
NAND2_X1 \myexu/_2925_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_2469_ ), .ZN(\myexu/_1944_ ) );
NAND2_X1 \myexu/_2926_ ( .A1(fanout_net_8 ), .A2(\myexu/_0305_ ), .ZN(\myexu/_1945_ ) );
NAND2_X1 \myexu/_2927_ ( .A1(\myexu/_1944_ ), .A2(\myexu/_1945_ ), .ZN(\myexu/_0012_ ) );
NAND2_X1 \myexu/_2928_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_2471_ ), .ZN(\myexu/_1946_ ) );
NAND2_X1 \myexu/_2929_ ( .A1(fanout_net_8 ), .A2(\myexu/_0307_ ), .ZN(\myexu/_1947_ ) );
NAND2_X1 \myexu/_2930_ ( .A1(\myexu/_1946_ ), .A2(\myexu/_1947_ ), .ZN(\myexu/_0014_ ) );
NOR2_X1 \myexu/_2931_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_0308_ ), .ZN(\myexu/_1948_ ) );
NOR2_X1 \myexu/_2932_ ( .A1(fanout_net_8 ), .A2(\myexu/_2472_ ), .ZN(\myexu/_1949_ ) );
NOR2_X1 \myexu/_2933_ ( .A1(\myexu/_1948_ ), .A2(\myexu/_1949_ ), .ZN(\myexu/_0015_ ) );
MUX2_X1 \myexu/_2934_ ( .A(\myexu/_2473_ ), .B(\myexu/_0309_ ), .S(fanout_net_8 ), .Z(\myexu/_0016_ ) );
NAND2_X1 \myexu/_2935_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_2474_ ), .ZN(\myexu/_1950_ ) );
NAND2_X1 \myexu/_2936_ ( .A1(fanout_net_8 ), .A2(\myexu/_0310_ ), .ZN(\myexu/_1951_ ) );
NAND2_X1 \myexu/_2937_ ( .A1(\myexu/_1950_ ), .A2(\myexu/_1951_ ), .ZN(\myexu/_0017_ ) );
MUX2_X1 \myexu/_2938_ ( .A(\myexu/_2475_ ), .B(\myexu/_0311_ ), .S(fanout_net_8 ), .Z(\myexu/_0018_ ) );
MUX2_X1 \myexu/_2939_ ( .A(\myexu/_2476_ ), .B(\myexu/_0312_ ), .S(fanout_net_8 ), .Z(\myexu/_0019_ ) );
MUX2_X1 \myexu/_2940_ ( .A(\myexu/_2477_ ), .B(\myexu/_0313_ ), .S(fanout_net_8 ), .Z(\myexu/_0020_ ) );
NAND2_X1 \myexu/_2941_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_2478_ ), .ZN(\myexu/_1952_ ) );
NAND2_X1 \myexu/_2942_ ( .A1(fanout_net_8 ), .A2(\myexu/_0314_ ), .ZN(\myexu/_1953_ ) );
NAND2_X1 \myexu/_2943_ ( .A1(\myexu/_1952_ ), .A2(\myexu/_1953_ ), .ZN(\myexu/_0021_ ) );
MUX2_X1 \myexu/_2944_ ( .A(\myexu/_2479_ ), .B(\myexu/_0315_ ), .S(\myexu/_2527_ ), .Z(\myexu/_0022_ ) );
NOR2_X1 \myexu/_2945_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_0316_ ), .ZN(\myexu/_1954_ ) );
NOR2_X1 \myexu/_2946_ ( .A1(\myexu/_2527_ ), .A2(\myexu/_2480_ ), .ZN(\myexu/_1955_ ) );
NOR2_X1 \myexu/_2947_ ( .A1(\myexu/_1954_ ), .A2(\myexu/_1955_ ), .ZN(\myexu/_0023_ ) );
NAND2_X1 \myexu/_2948_ ( .A1(\myexu/_1939_ ), .A2(\myexu/_2482_ ), .ZN(\myexu/_1956_ ) );
NAND2_X1 \myexu/_2949_ ( .A1(\myexu/_2527_ ), .A2(\myexu/_0318_ ), .ZN(\myexu/_1957_ ) );
NAND2_X1 \myexu/_2950_ ( .A1(\myexu/_1956_ ), .A2(\myexu/_1957_ ), .ZN(\myexu/_0025_ ) );
AND2_X2 \myexu/_2951_ ( .A1(\myexu/_2529_ ), .A2(\myexu/_2530_ ), .ZN(\myexu/_1958_ ) );
INV_X1 \myexu/_2952_ ( .A(\myexu/_1958_ ), .ZN(\myexu/_1959_ ) );
BUF_X4 \myexu/_2953_ ( .A(\myexu/_1959_ ), .Z(\myexu/_1960_ ) );
BUF_X4 \myexu/_2954_ ( .A(\myexu/_1960_ ), .Z(\myexu/_1961_ ) );
INV_X1 \myexu/_2955_ ( .A(\myexu/_2528_ ), .ZN(\myexu/_1962_ ) );
BUF_X4 \myexu/_2956_ ( .A(\myexu/_1962_ ), .Z(\myexu/_1963_ ) );
NOR2_X1 \myexu/_2957_ ( .A1(\myexu/_2427_ ), .A2(\myexu/_0295_ ), .ZN(\myexu/_1964_ ) );
AND2_X1 \myexu/_2958_ ( .A1(\myexu/_2427_ ), .A2(\myexu/_0295_ ), .ZN(\myexu/_1965_ ) );
OAI22_X1 \myexu/_2959_ ( .A1(\myexu/_1961_ ), .A2(\myexu/_1963_ ), .B1(\myexu/_1964_ ), .B2(\myexu/_1965_ ), .ZN(\myexu/_1966_ ) );
AND2_X2 \myexu/_2960_ ( .A1(\myexu/_1958_ ), .A2(\myexu/_1962_ ), .ZN(\myexu/_1967_ ) );
BUF_X4 \myexu/_2961_ ( .A(\myexu/_1967_ ), .Z(\myexu/_1968_ ) );
MUX2_X1 \myexu/_2962_ ( .A(\myexu/_1966_ ), .B(\myexu/_0243_ ), .S(\myexu/_1968_ ), .Z(\myexu/_1969_ ) );
INV_X1 \myexu/_2963_ ( .A(\myexu/_2536_ ), .ZN(\myexu/_1970_ ) );
NOR2_X1 \myexu/_2964_ ( .A1(\myexu/_1970_ ), .A2(\myexu/_2537_ ), .ZN(\myexu/_1971_ ) );
INV_X2 \myexu/_2965_ ( .A(fanout_net_5 ), .ZN(\myexu/_1972_ ) );
AND2_X1 \myexu/_2966_ ( .A1(\myexu/_1971_ ), .A2(\myexu/_1972_ ), .ZN(\myexu/_1973_ ) );
BUF_X4 \myexu/_2967_ ( .A(\myexu/_1973_ ), .Z(\myexu/_1974_ ) );
BUF_X4 \myexu/_2968_ ( .A(\myexu/_1974_ ), .Z(\myexu/_1975_ ) );
BUF_X4 \myexu/_2969_ ( .A(\myexu/_1975_ ), .Z(\myexu/_1976_ ) );
MUX2_X1 \myexu/_2970_ ( .A(\myexu/_0255_ ), .B(\myexu/_1969_ ), .S(\myexu/_1976_ ), .Z(\myexu/_0066_ ) );
XOR2_X1 \myexu/_2971_ ( .A(\myexu/_2438_ ), .B(\myexu/_0306_ ), .Z(\myexu/_1977_ ) );
XOR2_X1 \myexu/_2972_ ( .A(\myexu/_1977_ ), .B(\myexu/_1965_ ), .Z(\myexu/_1978_ ) );
BUF_X2 \myexu/_2973_ ( .A(\myexu/_1961_ ), .Z(\myexu/_1979_ ) );
NAND3_X1 \myexu/_2974_ ( .A1(\myexu/_1978_ ), .A2(\myexu/_1976_ ), .A3(\myexu/_1979_ ), .ZN(\myexu/_1980_ ) );
BUF_X8 \myexu/_2975_ ( .A(\myexu/_1971_ ), .Z(\myexu/_1981_ ) );
INV_X2 \myexu/_2976_ ( .A(\myexu/_1981_ ), .ZN(\myexu/_1982_ ) );
BUF_X4 \myexu/_2977_ ( .A(\myexu/_1982_ ), .Z(\myexu/_1983_ ) );
OAI21_X1 \myexu/_2978_ ( .A(\myexu/_0266_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1984_ ) );
BUF_X4 \myexu/_2979_ ( .A(\myexu/_1968_ ), .Z(\myexu/_1985_ ) );
BUF_X4 \myexu/_2980_ ( .A(\myexu/_1972_ ), .Z(\myexu/_1986_ ) );
BUF_X4 \myexu/_2981_ ( .A(\myexu/_1981_ ), .Z(\myexu/_1987_ ) );
BUF_X4 \myexu/_2982_ ( .A(\myexu/_1987_ ), .Z(\myexu/_1988_ ) );
NAND4_X1 \myexu/_2983_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_1986_ ), .A3(\myexu/_0246_ ), .A4(\myexu/_1988_ ), .ZN(\myexu/_1989_ ) );
NAND3_X1 \myexu/_2984_ ( .A1(\myexu/_1980_ ), .A2(\myexu/_1984_ ), .A3(\myexu/_1989_ ), .ZN(\myexu/_0067_ ) );
NAND2_X1 \myexu/_2985_ ( .A1(\myexu/_1977_ ), .A2(\myexu/_1965_ ), .ZN(\myexu/_1990_ ) );
INV_X1 \myexu/_2986_ ( .A(\myexu/_2438_ ), .ZN(\myexu/_1991_ ) );
INV_X1 \myexu/_2987_ ( .A(\myexu/_0306_ ), .ZN(\myexu/_1992_ ) );
OAI21_X1 \myexu/_2988_ ( .A(\myexu/_1990_ ), .B1(\myexu/_1991_ ), .B2(\myexu/_1992_ ), .ZN(\myexu/_1993_ ) );
XOR2_X1 \myexu/_2989_ ( .A(\myexu/_2449_ ), .B(\myexu/_0317_ ), .Z(\myexu/_1994_ ) );
XOR2_X1 \myexu/_2990_ ( .A(\myexu/_1993_ ), .B(\myexu/_1994_ ), .Z(\myexu/_1995_ ) );
NAND3_X1 \myexu/_2991_ ( .A1(\myexu/_1995_ ), .A2(\myexu/_1976_ ), .A3(\myexu/_1979_ ), .ZN(\myexu/_1996_ ) );
OAI21_X1 \myexu/_2992_ ( .A(\myexu/_0277_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1997_ ) );
NAND4_X1 \myexu/_2993_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_1986_ ), .A3(\myexu/_0247_ ), .A4(\myexu/_1988_ ), .ZN(\myexu/_1998_ ) );
NAND3_X1 \myexu/_2994_ ( .A1(\myexu/_1996_ ), .A2(\myexu/_1997_ ), .A3(\myexu/_1998_ ), .ZN(\myexu/_0068_ ) );
BUF_X4 \myexu/_2995_ ( .A(\myexu/_1982_ ), .Z(\myexu/_1999_ ) );
OAI21_X1 \myexu/_2996_ ( .A(\myexu/_0280_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_2000_ ) );
BUF_X4 \myexu/_2997_ ( .A(\myexu/_1972_ ), .Z(\myexu/_2001_ ) );
BUF_X4 \myexu/_2998_ ( .A(\myexu/_1981_ ), .Z(\myexu/_2002_ ) );
BUF_X4 \myexu/_2999_ ( .A(\myexu/_2002_ ), .Z(\myexu/_2003_ ) );
NAND4_X1 \myexu/_3000_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_2001_ ), .A3(\myexu/_0248_ ), .A4(\myexu/_2003_ ), .ZN(\myexu/_2004_ ) );
NAND2_X1 \myexu/_3001_ ( .A1(\myexu/_1993_ ), .A2(\myexu/_1994_ ), .ZN(\myexu/_2005_ ) );
NAND2_X1 \myexu/_3002_ ( .A1(\myexu/_2449_ ), .A2(\myexu/_0317_ ), .ZN(\myexu/_2006_ ) );
NAND2_X1 \myexu/_3003_ ( .A1(\myexu/_2005_ ), .A2(\myexu/_2006_ ), .ZN(\myexu/_2007_ ) );
AND2_X1 \myexu/_3004_ ( .A1(\myexu/_2452_ ), .A2(\myexu/_0320_ ), .ZN(\myexu/_2008_ ) );
NOR2_X1 \myexu/_3005_ ( .A1(\myexu/_2452_ ), .A2(\myexu/_0320_ ), .ZN(\myexu/_2009_ ) );
NOR2_X1 \myexu/_3006_ ( .A1(\myexu/_2008_ ), .A2(\myexu/_2009_ ), .ZN(\myexu/_2010_ ) );
XNOR2_X1 \myexu/_3007_ ( .A(\myexu/_2007_ ), .B(\myexu/_2010_ ), .ZN(\myexu/_2011_ ) );
BUF_X4 \myexu/_3008_ ( .A(\myexu/_1974_ ), .Z(\myexu/_2012_ ) );
NAND2_X1 \myexu/_3009_ ( .A1(\myexu/_2012_ ), .A2(\myexu/_1979_ ), .ZN(\myexu/_2013_ ) );
OAI211_X2 \myexu/_3010_ ( .A(\myexu/_2000_ ), .B(\myexu/_2004_ ), .C1(\myexu/_2011_ ), .C2(\myexu/_2013_ ), .ZN(\myexu/_0069_ ) );
AOI21_X1 \myexu/_3011_ ( .A(\myexu/_2009_ ), .B1(\myexu/_2005_ ), .B2(\myexu/_2006_ ), .ZN(\myexu/_2014_ ) );
OR2_X1 \myexu/_3012_ ( .A1(\myexu/_2014_ ), .A2(\myexu/_2008_ ), .ZN(\myexu/_2015_ ) );
XOR2_X1 \myexu/_3013_ ( .A(\myexu/_2453_ ), .B(\myexu/_0321_ ), .Z(\myexu/_2016_ ) );
XOR2_X1 \myexu/_3014_ ( .A(\myexu/_2015_ ), .B(\myexu/_2016_ ), .Z(\myexu/_2017_ ) );
NAND3_X1 \myexu/_3015_ ( .A1(\myexu/_2017_ ), .A2(\myexu/_1976_ ), .A3(\myexu/_1979_ ), .ZN(\myexu/_2018_ ) );
OAI21_X1 \myexu/_3016_ ( .A(\myexu/_0281_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_2019_ ) );
NAND4_X1 \myexu/_3017_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_1986_ ), .A3(\myexu/_0249_ ), .A4(\myexu/_1988_ ), .ZN(\myexu/_2020_ ) );
NAND3_X1 \myexu/_3018_ ( .A1(\myexu/_2018_ ), .A2(\myexu/_2019_ ), .A3(\myexu/_2020_ ), .ZN(\myexu/_0070_ ) );
AND2_X1 \myexu/_3019_ ( .A1(\myexu/_2453_ ), .A2(\myexu/_0321_ ), .ZN(\myexu/_2021_ ) );
AOI21_X1 \myexu/_3020_ ( .A(\myexu/_2021_ ), .B1(\myexu/_2015_ ), .B2(\myexu/_2016_ ), .ZN(\myexu/_2022_ ) );
XOR2_X1 \myexu/_3021_ ( .A(\myexu/_2454_ ), .B(\myexu/_0322_ ), .Z(\myexu/_2023_ ) );
XNOR2_X1 \myexu/_3022_ ( .A(\myexu/_2022_ ), .B(\myexu/_2023_ ), .ZN(\myexu/_2024_ ) );
NAND3_X1 \myexu/_3023_ ( .A1(\myexu/_2024_ ), .A2(\myexu/_1976_ ), .A3(\myexu/_1979_ ), .ZN(\myexu/_2025_ ) );
OAI21_X1 \myexu/_3024_ ( .A(\myexu/_0282_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_2026_ ) );
NAND4_X1 \myexu/_3025_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_1986_ ), .A3(\myexu/_0250_ ), .A4(\myexu/_1988_ ), .ZN(\myexu/_2027_ ) );
NAND3_X1 \myexu/_3026_ ( .A1(\myexu/_2025_ ), .A2(\myexu/_2026_ ), .A3(\myexu/_2027_ ), .ZN(\myexu/_0071_ ) );
AND2_X2 \myexu/_3027_ ( .A1(\myexu/_1958_ ), .A2(\myexu/_2528_ ), .ZN(\myexu/_2028_ ) );
INV_X2 \myexu/_3028_ ( .A(\myexu/_2028_ ), .ZN(\myexu/_2029_ ) );
BUF_X4 \myexu/_3029_ ( .A(\myexu/_2029_ ), .Z(\myexu/_2030_ ) );
BUF_X4 \myexu/_3030_ ( .A(\myexu/_2030_ ), .Z(\myexu/_2031_ ) );
BUF_X2 \myexu/_3031_ ( .A(\myexu/_1958_ ), .Z(\myexu/_2032_ ) );
BUF_X2 \myexu/_3032_ ( .A(\myexu/_2032_ ), .Z(\myexu/_2033_ ) );
BUF_X2 \myexu/_3033_ ( .A(\myexu/_1962_ ), .Z(\myexu/_2034_ ) );
NAND3_X1 \myexu/_3034_ ( .A1(\myexu/_2033_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_0251_ ), .ZN(\myexu/_2035_ ) );
NAND3_X1 \myexu/_3035_ ( .A1(\myexu/_2031_ ), .A2(\myexu/_2012_ ), .A3(\myexu/_2035_ ), .ZN(\myexu/_2036_ ) );
AND3_X1 \myexu/_3036_ ( .A1(\myexu/_2015_ ), .A2(\myexu/_2016_ ), .A3(\myexu/_2023_ ), .ZN(\myexu/_2037_ ) );
AND2_X1 \myexu/_3037_ ( .A1(\myexu/_2023_ ), .A2(\myexu/_2021_ ), .ZN(\myexu/_2038_ ) );
AOI21_X1 \myexu/_3038_ ( .A(\myexu/_2038_ ), .B1(\myexu/_2454_ ), .B2(\myexu/_0322_ ), .ZN(\myexu/_2039_ ) );
INV_X1 \myexu/_3039_ ( .A(\myexu/_2039_ ), .ZN(\myexu/_2040_ ) );
NOR2_X1 \myexu/_3040_ ( .A1(\myexu/_2037_ ), .A2(\myexu/_2040_ ), .ZN(\myexu/_2041_ ) );
XOR2_X1 \myexu/_3041_ ( .A(\myexu/_2455_ ), .B(\myexu/_0323_ ), .Z(\myexu/_2042_ ) );
XNOR2_X1 \myexu/_3042_ ( .A(\myexu/_2041_ ), .B(\myexu/_2042_ ), .ZN(\myexu/_2043_ ) );
AOI21_X1 \myexu/_3043_ ( .A(\myexu/_2036_ ), .B1(\myexu/_2043_ ), .B2(\myexu/_1979_ ), .ZN(\myexu/_2044_ ) );
BUF_X4 \myexu/_3044_ ( .A(\myexu/_1987_ ), .Z(\myexu/_2045_ ) );
CLKBUF_X2 \myexu/_3045_ ( .A(\myexu/_1972_ ), .Z(\myexu/_2046_ ) );
AOI21_X1 \myexu/_3046_ ( .A(\myexu/_0283_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_2046_ ), .ZN(\myexu/_2047_ ) );
NOR2_X1 \myexu/_3047_ ( .A1(\myexu/_2044_ ), .A2(\myexu/_2047_ ), .ZN(\myexu/_0072_ ) );
OAI21_X1 \myexu/_3048_ ( .A(\myexu/_0284_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_2048_ ) );
BUF_X4 \myexu/_3049_ ( .A(\myexu/_1967_ ), .Z(\myexu/_2049_ ) );
NAND4_X1 \myexu/_3050_ ( .A1(\myexu/_2049_ ), .A2(\myexu/_2001_ ), .A3(\myexu/_0252_ ), .A4(\myexu/_2003_ ), .ZN(\myexu/_2050_ ) );
NOR2_X1 \myexu/_3051_ ( .A1(\myexu/_2455_ ), .A2(\myexu/_0323_ ), .ZN(\myexu/_2051_ ) );
AND2_X1 \myexu/_3052_ ( .A1(\myexu/_2455_ ), .A2(\myexu/_0323_ ), .ZN(\myexu/_2052_ ) );
NOR3_X1 \myexu/_3053_ ( .A1(\myexu/_2041_ ), .A2(\myexu/_2051_ ), .A3(\myexu/_2052_ ), .ZN(\myexu/_2053_ ) );
OR2_X1 \myexu/_3054_ ( .A1(\myexu/_2053_ ), .A2(\myexu/_2052_ ), .ZN(\myexu/_2054_ ) );
XOR2_X1 \myexu/_3055_ ( .A(\myexu/_2456_ ), .B(\myexu/_0324_ ), .Z(\myexu/_2055_ ) );
XNOR2_X1 \myexu/_3056_ ( .A(\myexu/_2054_ ), .B(\myexu/_2055_ ), .ZN(\myexu/_2056_ ) );
OAI211_X2 \myexu/_3057_ ( .A(\myexu/_2048_ ), .B(\myexu/_2050_ ), .C1(\myexu/_2056_ ), .C2(\myexu/_2013_ ), .ZN(\myexu/_0073_ ) );
BUF_X4 \myexu/_3058_ ( .A(\myexu/_1958_ ), .Z(\myexu/_2057_ ) );
BUF_X4 \myexu/_3059_ ( .A(\myexu/_2057_ ), .Z(\myexu/_2058_ ) );
NAND3_X1 \myexu/_3060_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_0253_ ), .ZN(\myexu/_2059_ ) );
NAND3_X1 \myexu/_3061_ ( .A1(\myexu/_2031_ ), .A2(\myexu/_2012_ ), .A3(\myexu/_2059_ ), .ZN(\myexu/_2060_ ) );
AND2_X1 \myexu/_3062_ ( .A1(\myexu/_2042_ ), .A2(\myexu/_2055_ ), .ZN(\myexu/_2061_ ) );
OAI21_X1 \myexu/_3063_ ( .A(\myexu/_2061_ ), .B1(\myexu/_2037_ ), .B2(\myexu/_2040_ ), .ZN(\myexu/_2062_ ) );
AND2_X1 \myexu/_3064_ ( .A1(\myexu/_2055_ ), .A2(\myexu/_2052_ ), .ZN(\myexu/_2063_ ) );
AOI21_X1 \myexu/_3065_ ( .A(\myexu/_2063_ ), .B1(\myexu/_2456_ ), .B2(\myexu/_0324_ ), .ZN(\myexu/_2064_ ) );
AND2_X1 \myexu/_3066_ ( .A1(\myexu/_2062_ ), .A2(\myexu/_2064_ ), .ZN(\myexu/_2065_ ) );
XOR2_X1 \myexu/_3067_ ( .A(\myexu/_2457_ ), .B(\myexu/_0325_ ), .Z(\myexu/_2066_ ) );
XNOR2_X1 \myexu/_3068_ ( .A(\myexu/_2065_ ), .B(\myexu/_2066_ ), .ZN(\myexu/_2067_ ) );
AOI21_X1 \myexu/_3069_ ( .A(\myexu/_2060_ ), .B1(\myexu/_2067_ ), .B2(\myexu/_1979_ ), .ZN(\myexu/_2068_ ) );
AOI21_X1 \myexu/_3070_ ( .A(\myexu/_0285_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_2046_ ), .ZN(\myexu/_2069_ ) );
NOR2_X1 \myexu/_3071_ ( .A1(\myexu/_2068_ ), .A2(\myexu/_2069_ ), .ZN(\myexu/_0074_ ) );
BUF_X4 \myexu/_3072_ ( .A(\myexu/_2028_ ), .Z(\myexu/_2070_ ) );
INV_X1 \myexu/_3073_ ( .A(\myexu/_1974_ ), .ZN(\myexu/_2071_ ) );
BUF_X4 \myexu/_3074_ ( .A(\myexu/_2071_ ), .Z(\myexu/_2072_ ) );
AOI211_X4 \myexu/_3075_ ( .A(\myexu/_2070_ ), .B(\myexu/_2072_ ), .C1(\myexu/_0254_ ), .C2(\myexu/_1967_ ), .ZN(\myexu/_2073_ ) );
INV_X1 \myexu/_3076_ ( .A(\myexu/_2066_ ), .ZN(\myexu/_2074_ ) );
AOI21_X1 \myexu/_3077_ ( .A(\myexu/_2074_ ), .B1(\myexu/_2062_ ), .B2(\myexu/_2064_ ), .ZN(\myexu/_2075_ ) );
AND2_X1 \myexu/_3078_ ( .A1(\myexu/_2457_ ), .A2(\myexu/_0325_ ), .ZN(\myexu/_2076_ ) );
NOR2_X1 \myexu/_3079_ ( .A1(\myexu/_2075_ ), .A2(\myexu/_2076_ ), .ZN(\myexu/_2077_ ) );
XNOR2_X1 \myexu/_3080_ ( .A(\myexu/_2458_ ), .B(\myexu/_0326_ ), .ZN(\myexu/_2078_ ) );
XNOR2_X1 \myexu/_3081_ ( .A(\myexu/_2077_ ), .B(\myexu/_2078_ ), .ZN(\myexu/_2079_ ) );
BUF_X4 \myexu/_3082_ ( .A(\myexu/_2057_ ), .Z(\myexu/_2080_ ) );
OAI21_X1 \myexu/_3083_ ( .A(\myexu/_2073_ ), .B1(\myexu/_2079_ ), .B2(\myexu/_2080_ ), .ZN(\myexu/_2081_ ) );
CLKBUF_X2 \myexu/_3084_ ( .A(\myexu/_1974_ ), .Z(\myexu/_2082_ ) );
OR2_X1 \myexu/_3085_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_0286_ ), .ZN(\myexu/_2083_ ) );
AND2_X1 \myexu/_3086_ ( .A1(\myexu/_2081_ ), .A2(\myexu/_2083_ ), .ZN(\myexu/_0075_ ) );
AOI211_X4 \myexu/_3087_ ( .A(\myexu/_2074_ ), .B(\myexu/_2078_ ), .C1(\myexu/_2062_ ), .C2(\myexu/_2064_ ), .ZN(\myexu/_2084_ ) );
XOR2_X1 \myexu/_3088_ ( .A(\myexu/_2428_ ), .B(\myexu/_0296_ ), .Z(\myexu/_2085_ ) );
INV_X1 \myexu/_3089_ ( .A(\myexu/_2076_ ), .ZN(\myexu/_2086_ ) );
NOR2_X1 \myexu/_3090_ ( .A1(\myexu/_2078_ ), .A2(\myexu/_2086_ ), .ZN(\myexu/_2087_ ) );
AOI21_X1 \myexu/_3091_ ( .A(\myexu/_2087_ ), .B1(\myexu/_2458_ ), .B2(\myexu/_0326_ ), .ZN(\myexu/_2088_ ) );
INV_X1 \myexu/_3092_ ( .A(\myexu/_2088_ ), .ZN(\myexu/_2089_ ) );
OR3_X1 \myexu/_3093_ ( .A1(\myexu/_2084_ ), .A2(\myexu/_2085_ ), .A3(\myexu/_2089_ ), .ZN(\myexu/_2090_ ) );
OAI21_X1 \myexu/_3094_ ( .A(\myexu/_2085_ ), .B1(\myexu/_2084_ ), .B2(\myexu/_2089_ ), .ZN(\myexu/_2091_ ) );
NAND4_X1 \myexu/_3095_ ( .A1(\myexu/_2090_ ), .A2(\myexu/_1976_ ), .A3(\myexu/_1979_ ), .A4(\myexu/_2091_ ), .ZN(\myexu/_2092_ ) );
OAI21_X1 \myexu/_3096_ ( .A(\myexu/_0256_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_2093_ ) );
NAND4_X1 \myexu/_3097_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_1986_ ), .A3(\myexu/_0244_ ), .A4(\myexu/_1988_ ), .ZN(\myexu/_2094_ ) );
NAND3_X1 \myexu/_3098_ ( .A1(\myexu/_2092_ ), .A2(\myexu/_2093_ ), .A3(\myexu/_2094_ ), .ZN(\myexu/_0076_ ) );
OAI21_X1 \myexu/_3099_ ( .A(\myexu/_0257_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_2095_ ) );
NAND4_X1 \myexu/_3100_ ( .A1(\myexu/_2049_ ), .A2(\myexu/_2001_ ), .A3(\myexu/_0245_ ), .A4(\myexu/_2003_ ), .ZN(\myexu/_2096_ ) );
AND2_X1 \myexu/_3101_ ( .A1(\myexu/_2428_ ), .A2(\myexu/_0296_ ), .ZN(\myexu/_2097_ ) );
INV_X1 \myexu/_3102_ ( .A(\myexu/_2097_ ), .ZN(\myexu/_2098_ ) );
NAND2_X1 \myexu/_3103_ ( .A1(\myexu/_2091_ ), .A2(\myexu/_2098_ ), .ZN(\myexu/_2099_ ) );
XOR2_X1 \myexu/_3104_ ( .A(\myexu/_2429_ ), .B(\myexu/_0297_ ), .Z(\myexu/_2100_ ) );
XNOR2_X1 \myexu/_3105_ ( .A(\myexu/_2099_ ), .B(\myexu/_2100_ ), .ZN(\myexu/_2101_ ) );
OAI211_X2 \myexu/_3106_ ( .A(\myexu/_2095_ ), .B(\myexu/_2096_ ), .C1(\myexu/_2101_ ), .C2(\myexu/_2013_ ), .ZN(\myexu/_0077_ ) );
AOI21_X1 \myexu/_3107_ ( .A(\myexu/_2362_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_1986_ ), .ZN(\myexu/_2102_ ) );
INV_X1 \myexu/_3108_ ( .A(\myexu/_2459_ ), .ZN(\myexu/_2103_ ) );
BUF_X4 \myexu/_3109_ ( .A(\myexu/_2029_ ), .Z(\myexu/_2104_ ) );
INV_X1 \myexu/_3110_ ( .A(\myexu/_2260_ ), .ZN(\myexu/_2105_ ) );
OAI221_X1 \myexu/_3111_ ( .A(\myexu/_1975_ ), .B1(\myexu/_2103_ ), .B2(\myexu/_2057_ ), .C1(\myexu/_2104_ ), .C2(\myexu/_2105_ ), .ZN(\myexu/_2106_ ) );
INV_X1 \myexu/_3112_ ( .A(\myexu/_2524_ ), .ZN(\myexu/_2107_ ) );
NOR2_X1 \myexu/_3113_ ( .A1(\myexu/_2107_ ), .A2(\myexu/_2525_ ), .ZN(\myexu/_2108_ ) );
BUF_X4 \myexu/_3114_ ( .A(\myexu/_2108_ ), .Z(\myexu/_2109_ ) );
AND3_X1 \myexu/_3115_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1963_ ), .A3(\myexu/_2491_ ), .ZN(\myexu/_2110_ ) );
AOI21_X1 \myexu/_3116_ ( .A(\myexu/_2106_ ), .B1(\myexu/_2109_ ), .B2(\myexu/_2110_ ), .ZN(\myexu/_2111_ ) );
INV_X1 \myexu/_3117_ ( .A(\myexu/_2525_ ), .ZN(\myexu/_2112_ ) );
BUF_X2 \myexu/_3118_ ( .A(\myexu/_2112_ ), .Z(\myexu/_2113_ ) );
BUF_X4 \myexu/_3119_ ( .A(\myexu/_2113_ ), .Z(\myexu/_2114_ ) );
BUF_X4 \myexu/_3120_ ( .A(\myexu/_2114_ ), .Z(\myexu/_2115_ ) );
OAI211_X2 \myexu/_3121_ ( .A(\myexu/_2057_ ), .B(\myexu/_1963_ ), .C1(\myexu/_2115_ ), .C2(\myexu/_2491_ ), .ZN(\myexu/_2116_ ) );
NOR2_X1 \myexu/_3122_ ( .A1(\myexu/_2427_ ), .A2(fanout_net_7 ), .ZN(\myexu/_2117_ ) );
INV_X1 \myexu/_3123_ ( .A(fanout_net_7 ), .ZN(\myexu/_2118_ ) );
BUF_X4 \myexu/_3124_ ( .A(\myexu/_2118_ ), .Z(\myexu/_2119_ ) );
BUF_X4 \myexu/_3125_ ( .A(\myexu/_2119_ ), .Z(\myexu/_2120_ ) );
BUF_X4 \myexu/_3126_ ( .A(\myexu/_2120_ ), .Z(\myexu/_2121_ ) );
NOR2_X1 \myexu/_3127_ ( .A1(\myexu/_2121_ ), .A2(\myexu/_0295_ ), .ZN(\myexu/_2122_ ) );
OR3_X1 \myexu/_3128_ ( .A1(\myexu/_2116_ ), .A2(\myexu/_2117_ ), .A3(\myexu/_2122_ ), .ZN(\myexu/_2123_ ) );
AOI21_X1 \myexu/_3129_ ( .A(\myexu/_2102_ ), .B1(\myexu/_2111_ ), .B2(\myexu/_2123_ ), .ZN(\myexu/_0078_ ) );
AOI21_X1 \myexu/_3130_ ( .A(\myexu/_2373_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_1986_ ), .ZN(\myexu/_2124_ ) );
INV_X1 \myexu/_3131_ ( .A(\myexu/_2470_ ), .ZN(\myexu/_2125_ ) );
OAI211_X2 \myexu/_3132_ ( .A(\myexu/_1981_ ), .B(\myexu/_1972_ ), .C1(\myexu/_2032_ ), .C2(\myexu/_2125_ ), .ZN(\myexu/_2126_ ) );
BUF_X4 \myexu/_3133_ ( .A(\myexu/_2119_ ), .Z(\myexu/_2127_ ) );
NAND2_X1 \myexu/_3134_ ( .A1(\myexu/_1991_ ), .A2(\myexu/_2127_ ), .ZN(\myexu/_2128_ ) );
OAI221_X1 \myexu/_3135_ ( .A(\myexu/_2128_ ), .B1(\myexu/_0306_ ), .B2(\myexu/_2127_ ), .C1(\myexu/_2113_ ), .C2(\myexu/_2502_ ), .ZN(\myexu/_2129_ ) );
INV_X1 \myexu/_3136_ ( .A(\myexu/_1967_ ), .ZN(\myexu/_2130_ ) );
BUF_X4 \myexu/_3137_ ( .A(\myexu/_2130_ ), .Z(\myexu/_2131_ ) );
NOR2_X1 \myexu/_3138_ ( .A1(\myexu/_2129_ ), .A2(\myexu/_2131_ ), .ZN(\myexu/_2132_ ) );
BUF_X4 \myexu/_3139_ ( .A(\myexu/_2028_ ), .Z(\myexu/_2133_ ) );
AOI211_X4 \myexu/_3140_ ( .A(\myexu/_2126_ ), .B(\myexu/_2132_ ), .C1(\myexu/_2271_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_2134_ ) );
NAND3_X1 \myexu/_3141_ ( .A1(\myexu/_1985_ ), .A2(\myexu/_2502_ ), .A3(\myexu/_2109_ ), .ZN(\myexu/_2135_ ) );
AOI21_X1 \myexu/_3142_ ( .A(\myexu/_2124_ ), .B1(\myexu/_2134_ ), .B2(\myexu/_2135_ ), .ZN(\myexu/_0079_ ) );
AOI221_X4 \myexu/_3143_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2481_ ), .B2(\myexu/_1961_ ), .C1(\myexu/_2282_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_2136_ ) );
INV_X1 \myexu/_3144_ ( .A(\myexu/_2449_ ), .ZN(\myexu/_2137_ ) );
NAND2_X1 \myexu/_3145_ ( .A1(\myexu/_2137_ ), .A2(\myexu/_2121_ ), .ZN(\myexu/_2138_ ) );
OAI221_X1 \myexu/_3146_ ( .A(\myexu/_2138_ ), .B1(\myexu/_0317_ ), .B2(\myexu/_2121_ ), .C1(\myexu/_2114_ ), .C2(\myexu/_2513_ ), .ZN(\myexu/_2139_ ) );
BUF_X2 \myexu/_3147_ ( .A(\myexu/_2130_ ), .Z(\myexu/_2140_ ) );
OR2_X1 \myexu/_3148_ ( .A1(\myexu/_2139_ ), .A2(\myexu/_2140_ ), .ZN(\myexu/_2141_ ) );
NAND3_X1 \myexu/_3149_ ( .A1(\myexu/_2049_ ), .A2(\myexu/_2513_ ), .A3(\myexu/_2109_ ), .ZN(\myexu/_2142_ ) );
NAND3_X1 \myexu/_3150_ ( .A1(\myexu/_2136_ ), .A2(\myexu/_2141_ ), .A3(\myexu/_2142_ ), .ZN(\myexu/_2143_ ) );
OR2_X1 \myexu/_3151_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2384_ ), .ZN(\myexu/_2144_ ) );
AND2_X1 \myexu/_3152_ ( .A1(\myexu/_2143_ ), .A2(\myexu/_2144_ ), .ZN(\myexu/_0080_ ) );
NOR2_X1 \myexu/_3153_ ( .A1(\myexu/_2452_ ), .A2(fanout_net_7 ), .ZN(\myexu/_2145_ ) );
INV_X1 \myexu/_3154_ ( .A(\myexu/_2516_ ), .ZN(\myexu/_2146_ ) );
AOI221_X4 \myexu/_3155_ ( .A(\myexu/_2145_ ), .B1(\myexu/_1931_ ), .B2(fanout_net_7 ), .C1(\myexu/_2525_ ), .C2(\myexu/_2146_ ), .ZN(\myexu/_2147_ ) );
AND3_X1 \myexu/_3156_ ( .A1(\myexu/_2113_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2516_ ), .ZN(\myexu/_2148_ ) );
OAI21_X1 \myexu/_3157_ ( .A(\myexu/_1968_ ), .B1(\myexu/_2147_ ), .B2(\myexu/_2148_ ), .ZN(\myexu/_2149_ ) );
INV_X1 \myexu/_3158_ ( .A(\myexu/_2285_ ), .ZN(\myexu/_2150_ ) );
OAI221_X1 \myexu/_3159_ ( .A(\myexu/_2149_ ), .B1(\myexu/_1929_ ), .B2(\myexu/_2058_ ), .C1(\myexu/_2150_ ), .C2(\myexu/_2104_ ), .ZN(\myexu/_2151_ ) );
MUX2_X1 \myexu/_3160_ ( .A(\myexu/_2387_ ), .B(\myexu/_2151_ ), .S(\myexu/_1976_ ), .Z(\myexu/_0081_ ) );
AOI221_X4 \myexu/_3161_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2485_ ), .B2(\myexu/_1961_ ), .C1(\myexu/_2286_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_2152_ ) );
CLKBUF_X2 \myexu/_3162_ ( .A(\myexu/_2120_ ), .Z(\myexu/_2153_ ) );
OR2_X1 \myexu/_3163_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0321_ ), .ZN(\myexu/_2154_ ) );
OAI221_X1 \myexu/_3164_ ( .A(\myexu/_2154_ ), .B1(\myexu/_2453_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2517_ ), .ZN(\myexu/_2155_ ) );
CLKBUF_X2 \myexu/_3165_ ( .A(\myexu/_2130_ ), .Z(\myexu/_2156_ ) );
OR2_X1 \myexu/_3166_ ( .A1(\myexu/_2155_ ), .A2(\myexu/_2156_ ), .ZN(\myexu/_2157_ ) );
BUF_X2 \myexu/_3167_ ( .A(\myexu/_1967_ ), .Z(\myexu/_2158_ ) );
NAND3_X1 \myexu/_3168_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2517_ ), .A3(\myexu/_2109_ ), .ZN(\myexu/_2159_ ) );
NAND3_X1 \myexu/_3169_ ( .A1(\myexu/_2152_ ), .A2(\myexu/_2157_ ), .A3(\myexu/_2159_ ), .ZN(\myexu/_2160_ ) );
OR2_X1 \myexu/_3170_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2388_ ), .ZN(\myexu/_2161_ ) );
AND2_X1 \myexu/_3171_ ( .A1(\myexu/_2160_ ), .A2(\myexu/_2161_ ), .ZN(\myexu/_0082_ ) );
AOI221_X4 \myexu/_3172_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2486_ ), .B2(\myexu/_1961_ ), .C1(\myexu/_2287_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_2162_ ) );
NAND3_X1 \myexu/_3173_ ( .A1(\myexu/_2049_ ), .A2(\myexu/_2518_ ), .A3(\myexu/_2109_ ), .ZN(\myexu/_2163_ ) );
INV_X1 \myexu/_3174_ ( .A(\myexu/_0322_ ), .ZN(\myexu/_2164_ ) );
NAND2_X1 \myexu/_3175_ ( .A1(\myexu/_2164_ ), .A2(fanout_net_7 ), .ZN(\myexu/_2165_ ) );
OAI221_X1 \myexu/_3176_ ( .A(\myexu/_2165_ ), .B1(\myexu/_2454_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2518_ ), .ZN(\myexu/_2166_ ) );
OR2_X1 \myexu/_3177_ ( .A1(\myexu/_2140_ ), .A2(\myexu/_2166_ ), .ZN(\myexu/_2167_ ) );
NAND3_X1 \myexu/_3178_ ( .A1(\myexu/_2162_ ), .A2(\myexu/_2163_ ), .A3(\myexu/_2167_ ), .ZN(\myexu/_2168_ ) );
OR2_X1 \myexu/_3179_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2389_ ), .ZN(\myexu/_2169_ ) );
AND2_X1 \myexu/_3180_ ( .A1(\myexu/_2168_ ), .A2(\myexu/_2169_ ), .ZN(\myexu/_0083_ ) );
NOR2_X1 \myexu/_3181_ ( .A1(\myexu/_2119_ ), .A2(\myexu/_0323_ ), .ZN(\myexu/_2170_ ) );
INV_X1 \myexu/_3182_ ( .A(\myexu/_2455_ ), .ZN(\myexu/_2171_ ) );
INV_X1 \myexu/_3183_ ( .A(\myexu/_2519_ ), .ZN(\myexu/_2172_ ) );
AOI221_X4 \myexu/_3184_ ( .A(\myexu/_2170_ ), .B1(\myexu/_2171_ ), .B2(\myexu/_2120_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_2172_ ), .ZN(\myexu/_2173_ ) );
AND3_X1 \myexu/_3185_ ( .A1(\myexu/_2113_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2519_ ), .ZN(\myexu/_2174_ ) );
OAI21_X1 \myexu/_3186_ ( .A(\myexu/_1968_ ), .B1(\myexu/_2173_ ), .B2(\myexu/_2174_ ), .ZN(\myexu/_2175_ ) );
INV_X1 \myexu/_3187_ ( .A(\myexu/_2487_ ), .ZN(\myexu/_2176_ ) );
INV_X1 \myexu/_3188_ ( .A(\myexu/_2288_ ), .ZN(\myexu/_2177_ ) );
OAI221_X1 \myexu/_3189_ ( .A(\myexu/_2175_ ), .B1(\myexu/_2176_ ), .B2(\myexu/_2057_ ), .C1(\myexu/_2177_ ), .C2(\myexu/_2104_ ), .ZN(\myexu/_2178_ ) );
MUX2_X1 \myexu/_3190_ ( .A(\myexu/_2390_ ), .B(\myexu/_2178_ ), .S(\myexu/_1976_ ), .Z(\myexu/_0084_ ) );
AOI221_X4 \myexu/_3191_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2488_ ), .B2(\myexu/_1961_ ), .C1(\myexu/_2289_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_2179_ ) );
NOR2_X1 \myexu/_3192_ ( .A1(\myexu/_2127_ ), .A2(\myexu/_0324_ ), .ZN(\myexu/_2180_ ) );
INV_X1 \myexu/_3193_ ( .A(\myexu/_2456_ ), .ZN(\myexu/_2181_ ) );
INV_X1 \myexu/_3194_ ( .A(\myexu/_2520_ ), .ZN(\myexu/_2182_ ) );
AOI221_X4 \myexu/_3195_ ( .A(\myexu/_2180_ ), .B1(\myexu/_2181_ ), .B2(\myexu/_2127_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_2182_ ), .ZN(\myexu/_2183_ ) );
NAND2_X1 \myexu/_3196_ ( .A1(\myexu/_2183_ ), .A2(\myexu/_2049_ ), .ZN(\myexu/_2184_ ) );
NAND3_X1 \myexu/_3197_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2520_ ), .A3(\myexu/_2109_ ), .ZN(\myexu/_2185_ ) );
NAND3_X1 \myexu/_3198_ ( .A1(\myexu/_2179_ ), .A2(\myexu/_2184_ ), .A3(\myexu/_2185_ ), .ZN(\myexu/_2186_ ) );
OR2_X1 \myexu/_3199_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2391_ ), .ZN(\myexu/_2187_ ) );
AND2_X1 \myexu/_3200_ ( .A1(\myexu/_2186_ ), .A2(\myexu/_2187_ ), .ZN(\myexu/_0085_ ) );
AOI221_X4 \myexu/_3201_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2489_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2290_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_2188_ ) );
OR2_X1 \myexu/_3202_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0325_ ), .ZN(\myexu/_2189_ ) );
OAI221_X1 \myexu/_3203_ ( .A(\myexu/_2189_ ), .B1(\myexu/_2457_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2521_ ), .ZN(\myexu/_2190_ ) );
OR2_X1 \myexu/_3204_ ( .A1(\myexu/_2190_ ), .A2(\myexu/_2156_ ), .ZN(\myexu/_2191_ ) );
BUF_X2 \myexu/_3205_ ( .A(\myexu/_2108_ ), .Z(\myexu/_2192_ ) );
NAND3_X1 \myexu/_3206_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2521_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_2193_ ) );
NAND3_X1 \myexu/_3207_ ( .A1(\myexu/_2188_ ), .A2(\myexu/_2191_ ), .A3(\myexu/_2193_ ), .ZN(\myexu/_2194_ ) );
OR2_X1 \myexu/_3208_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2392_ ), .ZN(\myexu/_2195_ ) );
AND2_X1 \myexu/_3209_ ( .A1(\myexu/_2194_ ), .A2(\myexu/_2195_ ), .ZN(\myexu/_0086_ ) );
NOR2_X1 \myexu/_3210_ ( .A1(\myexu/_2119_ ), .A2(\myexu/_0326_ ), .ZN(\myexu/_2196_ ) );
INV_X1 \myexu/_3211_ ( .A(\myexu/_2458_ ), .ZN(\myexu/_2197_ ) );
INV_X1 \myexu/_3212_ ( .A(\myexu/_2522_ ), .ZN(\myexu/_2198_ ) );
AOI221_X4 \myexu/_3213_ ( .A(\myexu/_2196_ ), .B1(\myexu/_2197_ ), .B2(\myexu/_2120_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_2198_ ), .ZN(\myexu/_2199_ ) );
AND3_X1 \myexu/_3214_ ( .A1(\myexu/_2113_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2522_ ), .ZN(\myexu/_2200_ ) );
OAI21_X1 \myexu/_3215_ ( .A(\myexu/_1968_ ), .B1(\myexu/_2199_ ), .B2(\myexu/_2200_ ), .ZN(\myexu/_2201_ ) );
INV_X1 \myexu/_3216_ ( .A(\myexu/_2490_ ), .ZN(\myexu/_2202_ ) );
INV_X1 \myexu/_3217_ ( .A(\myexu/_2291_ ), .ZN(\myexu/_2203_ ) );
OAI221_X1 \myexu/_3218_ ( .A(\myexu/_2201_ ), .B1(\myexu/_2202_ ), .B2(\myexu/_2057_ ), .C1(\myexu/_2203_ ), .C2(\myexu/_2104_ ), .ZN(\myexu/_2204_ ) );
BUF_X4 \myexu/_3219_ ( .A(\myexu/_1975_ ), .Z(\myexu/_2205_ ) );
MUX2_X1 \myexu/_3220_ ( .A(\myexu/_2393_ ), .B(\myexu/_2204_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0087_ ) );
AOI21_X1 \myexu/_3221_ ( .A(\myexu/_2363_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_1986_ ), .ZN(\myexu/_2206_ ) );
CLKBUF_X2 \myexu/_3222_ ( .A(\myexu/_1960_ ), .Z(\myexu/_2207_ ) );
AOI221_X4 \myexu/_3223_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2460_ ), .B2(\myexu/_2207_ ), .C1(\myexu/_2261_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_2208_ ) );
NOR2_X1 \myexu/_3224_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0296_ ), .ZN(\myexu/_2209_ ) );
INV_X1 \myexu/_3225_ ( .A(\myexu/_2428_ ), .ZN(\myexu/_2210_ ) );
INV_X1 \myexu/_3226_ ( .A(\myexu/_2492_ ), .ZN(\myexu/_2211_ ) );
AOI221_X4 \myexu/_3227_ ( .A(\myexu/_2209_ ), .B1(\myexu/_2210_ ), .B2(\myexu/_2121_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_2211_ ), .ZN(\myexu/_2212_ ) );
AND3_X1 \myexu/_3228_ ( .A1(\myexu/_2115_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2492_ ), .ZN(\myexu/_2213_ ) );
OAI21_X1 \myexu/_3229_ ( .A(\myexu/_1985_ ), .B1(\myexu/_2212_ ), .B2(\myexu/_2213_ ), .ZN(\myexu/_2214_ ) );
AOI21_X1 \myexu/_3230_ ( .A(\myexu/_2206_ ), .B1(\myexu/_2208_ ), .B2(\myexu/_2214_ ), .ZN(\myexu/_0088_ ) );
AOI221_X4 \myexu/_3231_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2461_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2262_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_2215_ ) );
AND3_X1 \myexu/_3232_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1963_ ), .A3(\myexu/_2493_ ), .ZN(\myexu/_2216_ ) );
NAND2_X1 \myexu/_3233_ ( .A1(\myexu/_2216_ ), .A2(\myexu/_2109_ ), .ZN(\myexu/_2217_ ) );
OR2_X1 \myexu/_3234_ ( .A1(\myexu/_2127_ ), .A2(\myexu/_0297_ ), .ZN(\myexu/_2218_ ) );
OAI221_X1 \myexu/_3235_ ( .A(\myexu/_2218_ ), .B1(\myexu/_2429_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2493_ ), .ZN(\myexu/_2219_ ) );
OR2_X1 \myexu/_3236_ ( .A1(\myexu/_2219_ ), .A2(\myexu/_2156_ ), .ZN(\myexu/_2220_ ) );
NAND3_X1 \myexu/_3237_ ( .A1(\myexu/_2215_ ), .A2(\myexu/_2217_ ), .A3(\myexu/_2220_ ), .ZN(\myexu/_2221_ ) );
OR2_X1 \myexu/_3238_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2364_ ), .ZN(\myexu/_2222_ ) );
AND2_X1 \myexu/_3239_ ( .A1(\myexu/_2221_ ), .A2(\myexu/_2222_ ), .ZN(\myexu/_0089_ ) );
AOI21_X1 \myexu/_3240_ ( .A(\myexu/_2365_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_1986_ ), .ZN(\myexu/_2223_ ) );
AOI221_X4 \myexu/_3241_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2462_ ), .B2(\myexu/_2207_ ), .C1(\myexu/_2263_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_2224_ ) );
NOR2_X1 \myexu/_3242_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0298_ ), .ZN(\myexu/_2225_ ) );
INV_X1 \myexu/_3243_ ( .A(\myexu/_2430_ ), .ZN(\myexu/_2226_ ) );
INV_X1 \myexu/_3244_ ( .A(\myexu/_2494_ ), .ZN(\myexu/_2227_ ) );
AOI221_X4 \myexu/_3245_ ( .A(\myexu/_2225_ ), .B1(\myexu/_2226_ ), .B2(\myexu/_2153_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_2227_ ), .ZN(\myexu/_2228_ ) );
AND3_X1 \myexu/_3246_ ( .A1(\myexu/_2115_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2494_ ), .ZN(\myexu/_2229_ ) );
OAI21_X1 \myexu/_3247_ ( .A(\myexu/_1985_ ), .B1(\myexu/_2228_ ), .B2(\myexu/_2229_ ), .ZN(\myexu/_2230_ ) );
AOI21_X1 \myexu/_3248_ ( .A(\myexu/_2223_ ), .B1(\myexu/_2224_ ), .B2(\myexu/_2230_ ), .ZN(\myexu/_0090_ ) );
AOI21_X1 \myexu/_3249_ ( .A(\myexu/_2366_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_1986_ ), .ZN(\myexu/_2231_ ) );
AOI211_X4 \myexu/_3250_ ( .A(fanout_net_5 ), .B(\myexu/_1982_ ), .C1(\myexu/_2463_ ), .C2(\myexu/_1961_ ), .ZN(\myexu/_2232_ ) );
INV_X1 \myexu/_3251_ ( .A(\myexu/_2264_ ), .ZN(\myexu/_2233_ ) );
BUF_X4 \myexu/_3252_ ( .A(\myexu/_2029_ ), .Z(\myexu/_2234_ ) );
OAI21_X1 \myexu/_3253_ ( .A(\myexu/_2232_ ), .B1(\myexu/_2233_ ), .B2(\myexu/_2234_ ), .ZN(\myexu/_2235_ ) );
AND3_X1 \myexu/_3254_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1963_ ), .A3(\myexu/_2495_ ), .ZN(\myexu/_2236_ ) );
AOI21_X1 \myexu/_3255_ ( .A(\myexu/_2235_ ), .B1(\myexu/_2109_ ), .B2(\myexu/_2236_ ), .ZN(\myexu/_2237_ ) );
OAI211_X2 \myexu/_3256_ ( .A(\myexu/_2057_ ), .B(\myexu/_1963_ ), .C1(\myexu/_2115_ ), .C2(\myexu/_2495_ ), .ZN(\myexu/_2238_ ) );
NOR2_X1 \myexu/_3257_ ( .A1(\myexu/_2431_ ), .A2(fanout_net_7 ), .ZN(\myexu/_2239_ ) );
NOR2_X1 \myexu/_3258_ ( .A1(\myexu/_2121_ ), .A2(\myexu/_0299_ ), .ZN(\myexu/_2240_ ) );
OR3_X1 \myexu/_3259_ ( .A1(\myexu/_2238_ ), .A2(\myexu/_2239_ ), .A3(\myexu/_2240_ ), .ZN(\myexu/_2241_ ) );
AOI21_X1 \myexu/_3260_ ( .A(\myexu/_2231_ ), .B1(\myexu/_2237_ ), .B2(\myexu/_2241_ ), .ZN(\myexu/_0091_ ) );
AOI221_X4 \myexu/_3261_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2464_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2265_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_2242_ ) );
OR2_X1 \myexu/_3262_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0300_ ), .ZN(\myexu/_2243_ ) );
OAI221_X1 \myexu/_3263_ ( .A(\myexu/_2243_ ), .B1(\myexu/_2432_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2496_ ), .ZN(\myexu/_2244_ ) );
OR2_X1 \myexu/_3264_ ( .A1(\myexu/_2244_ ), .A2(\myexu/_2156_ ), .ZN(\myexu/_2245_ ) );
NAND3_X1 \myexu/_3265_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2496_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_2246_ ) );
NAND3_X1 \myexu/_3266_ ( .A1(\myexu/_2242_ ), .A2(\myexu/_2245_ ), .A3(\myexu/_2246_ ), .ZN(\myexu/_2247_ ) );
OR2_X1 \myexu/_3267_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2367_ ), .ZN(\myexu/_2248_ ) );
AND2_X1 \myexu/_3268_ ( .A1(\myexu/_2247_ ), .A2(\myexu/_2248_ ), .ZN(\myexu/_0092_ ) );
NOR2_X1 \myexu/_3269_ ( .A1(\myexu/_2433_ ), .A2(fanout_net_7 ), .ZN(\myexu/_2249_ ) );
NOR2_X1 \myexu/_3270_ ( .A1(\myexu/_2120_ ), .A2(\myexu/_0301_ ), .ZN(\myexu/_2250_ ) );
INV_X1 \myexu/_3271_ ( .A(\myexu/_2497_ ), .ZN(\myexu/_2251_ ) );
AOI211_X4 \myexu/_3272_ ( .A(\myexu/_2249_ ), .B(\myexu/_2250_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_2251_ ), .ZN(\myexu/_2252_ ) );
AND3_X1 \myexu/_3273_ ( .A1(\myexu/_2113_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2497_ ), .ZN(\myexu/_2253_ ) );
OAI21_X1 \myexu/_3274_ ( .A(\myexu/_1968_ ), .B1(\myexu/_2252_ ), .B2(\myexu/_2253_ ), .ZN(\myexu/_2254_ ) );
INV_X1 \myexu/_3275_ ( .A(\myexu/_2465_ ), .ZN(\myexu/_2255_ ) );
INV_X1 \myexu/_3276_ ( .A(\myexu/_2266_ ), .ZN(\myexu/_2256_ ) );
OAI221_X1 \myexu/_3277_ ( .A(\myexu/_2254_ ), .B1(\myexu/_2255_ ), .B2(\myexu/_2057_ ), .C1(\myexu/_2256_ ), .C2(\myexu/_2104_ ), .ZN(\myexu/_2257_ ) );
MUX2_X1 \myexu/_3278_ ( .A(\myexu/_2368_ ), .B(\myexu/_2257_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0093_ ) );
AOI221_X4 \myexu/_3279_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2466_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2267_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_2258_ ) );
OR2_X1 \myexu/_3280_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0302_ ), .ZN(\myexu/_2259_ ) );
OAI221_X1 \myexu/_3281_ ( .A(\myexu/_2259_ ), .B1(\myexu/_2434_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2498_ ), .ZN(\myexu/_0327_ ) );
OR2_X1 \myexu/_3282_ ( .A1(\myexu/_0327_ ), .A2(\myexu/_2156_ ), .ZN(\myexu/_0328_ ) );
NAND3_X1 \myexu/_3283_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2498_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_0329_ ) );
NAND3_X1 \myexu/_3284_ ( .A1(\myexu/_2258_ ), .A2(\myexu/_0328_ ), .A3(\myexu/_0329_ ), .ZN(\myexu/_0330_ ) );
OR2_X1 \myexu/_3285_ ( .A1(\myexu/_2082_ ), .A2(\myexu/_2369_ ), .ZN(\myexu/_0331_ ) );
AND2_X1 \myexu/_3286_ ( .A1(\myexu/_0330_ ), .A2(\myexu/_0331_ ), .ZN(\myexu/_0094_ ) );
AOI21_X1 \myexu/_3287_ ( .A(\myexu/_2370_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_2001_ ), .ZN(\myexu/_0332_ ) );
INV_X1 \myexu/_3288_ ( .A(\myexu/_2435_ ), .ZN(\myexu/_0333_ ) );
NAND2_X1 \myexu/_3289_ ( .A1(\myexu/_0333_ ), .A2(\myexu/_2127_ ), .ZN(\myexu/_0334_ ) );
OAI221_X1 \myexu/_3290_ ( .A(\myexu/_0334_ ), .B1(\myexu/_0303_ ), .B2(\myexu/_2127_ ), .C1(\myexu/_2113_ ), .C2(\myexu/_2499_ ), .ZN(\myexu/_0335_ ) );
NOR2_X1 \myexu/_3291_ ( .A1(\myexu/_0335_ ), .A2(\myexu/_2131_ ), .ZN(\myexu/_0336_ ) );
AOI221_X4 \myexu/_3292_ ( .A(\myexu/_0336_ ), .B1(\myexu/_2467_ ), .B2(\myexu/_2207_ ), .C1(\myexu/_2268_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_0337_ ) );
AND3_X1 \myexu/_3293_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1962_ ), .A3(\myexu/_2499_ ), .ZN(\myexu/_0338_ ) );
AOI211_X4 \myexu/_3294_ ( .A(fanout_net_5 ), .B(\myexu/_1982_ ), .C1(\myexu/_0338_ ), .C2(\myexu/_2108_ ), .ZN(\myexu/_0339_ ) );
AOI21_X1 \myexu/_3295_ ( .A(\myexu/_0332_ ), .B1(\myexu/_0337_ ), .B2(\myexu/_0339_ ), .ZN(\myexu/_0095_ ) );
AOI21_X1 \myexu/_3296_ ( .A(\myexu/_2371_ ), .B1(\myexu/_1988_ ), .B2(\myexu/_2001_ ), .ZN(\myexu/_0340_ ) );
AOI221_X4 \myexu/_3297_ ( .A(\myexu/_2072_ ), .B1(\myexu/_2468_ ), .B2(\myexu/_1961_ ), .C1(\myexu/_2269_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_0341_ ) );
INV_X1 \myexu/_3298_ ( .A(\myexu/_2436_ ), .ZN(\myexu/_0342_ ) );
NOR2_X1 \myexu/_3299_ ( .A1(\myexu/_0342_ ), .A2(fanout_net_7 ), .ZN(\myexu/_0343_ ) );
AOI221_X4 \myexu/_3300_ ( .A(\myexu/_0343_ ), .B1(\myexu/_0304_ ), .B2(fanout_net_7 ), .C1(\myexu/_2500_ ), .C2(\myexu/_2108_ ), .ZN(\myexu/_0344_ ) );
NOR2_X1 \myexu/_3301_ ( .A1(\myexu/_2115_ ), .A2(\myexu/_2500_ ), .ZN(\myexu/_0345_ ) );
OR3_X1 \myexu/_3302_ ( .A1(\myexu/_0344_ ), .A2(\myexu/_2140_ ), .A3(\myexu/_0345_ ), .ZN(\myexu/_0346_ ) );
AOI21_X1 \myexu/_3303_ ( .A(\myexu/_0340_ ), .B1(\myexu/_0341_ ), .B2(\myexu/_0346_ ), .ZN(\myexu/_0096_ ) );
NOR2_X1 \myexu/_3304_ ( .A1(\myexu/_2119_ ), .A2(\myexu/_0305_ ), .ZN(\myexu/_0347_ ) );
INV_X1 \myexu/_3305_ ( .A(\myexu/_2437_ ), .ZN(\myexu/_0348_ ) );
INV_X1 \myexu/_3306_ ( .A(\myexu/_2501_ ), .ZN(\myexu/_0349_ ) );
AOI221_X4 \myexu/_3307_ ( .A(\myexu/_0347_ ), .B1(\myexu/_0348_ ), .B2(\myexu/_2120_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0349_ ), .ZN(\myexu/_0350_ ) );
AND3_X1 \myexu/_3308_ ( .A1(\myexu/_2113_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2501_ ), .ZN(\myexu/_0351_ ) );
OAI21_X1 \myexu/_3309_ ( .A(\myexu/_1968_ ), .B1(\myexu/_0350_ ), .B2(\myexu/_0351_ ), .ZN(\myexu/_0352_ ) );
INV_X1 \myexu/_3310_ ( .A(\myexu/_2469_ ), .ZN(\myexu/_0353_ ) );
INV_X1 \myexu/_3311_ ( .A(\myexu/_2270_ ), .ZN(\myexu/_0354_ ) );
OAI221_X1 \myexu/_3312_ ( .A(\myexu/_0352_ ), .B1(\myexu/_0353_ ), .B2(\myexu/_2057_ ), .C1(\myexu/_0354_ ), .C2(\myexu/_2030_ ), .ZN(\myexu/_0355_ ) );
MUX2_X1 \myexu/_3313_ ( .A(\myexu/_2372_ ), .B(\myexu/_0355_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0097_ ) );
AOI221_X4 \myexu/_3314_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2471_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2272_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_0356_ ) );
OR2_X1 \myexu/_3315_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0307_ ), .ZN(\myexu/_0357_ ) );
OAI221_X1 \myexu/_3316_ ( .A(\myexu/_0357_ ), .B1(\myexu/_2439_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2503_ ), .ZN(\myexu/_0358_ ) );
OR2_X1 \myexu/_3317_ ( .A1(\myexu/_0358_ ), .A2(\myexu/_2156_ ), .ZN(\myexu/_0359_ ) );
NAND3_X1 \myexu/_3318_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2503_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_0360_ ) );
NAND3_X1 \myexu/_3319_ ( .A1(\myexu/_0356_ ), .A2(\myexu/_0359_ ), .A3(\myexu/_0360_ ), .ZN(\myexu/_0361_ ) );
OR2_X1 \myexu/_3320_ ( .A1(\myexu/_1975_ ), .A2(\myexu/_2374_ ), .ZN(\myexu/_0362_ ) );
AND2_X1 \myexu/_3321_ ( .A1(\myexu/_0361_ ), .A2(\myexu/_0362_ ), .ZN(\myexu/_0098_ ) );
INV_X1 \myexu/_3322_ ( .A(\myexu/_2472_ ), .ZN(\myexu/_0363_ ) );
INV_X1 \myexu/_3323_ ( .A(\myexu/_2273_ ), .ZN(\myexu/_0364_ ) );
OAI221_X1 \myexu/_3324_ ( .A(\myexu/_1974_ ), .B1(\myexu/_0363_ ), .B2(\myexu/_1958_ ), .C1(\myexu/_2029_ ), .C2(\myexu/_0364_ ), .ZN(\myexu/_0365_ ) );
NOR2_X1 \myexu/_3325_ ( .A1(\myexu/_2119_ ), .A2(\myexu/_0308_ ), .ZN(\myexu/_0366_ ) );
INV_X1 \myexu/_3326_ ( .A(\myexu/_2440_ ), .ZN(\myexu/_0367_ ) );
INV_X1 \myexu/_3327_ ( .A(\myexu/_2504_ ), .ZN(\myexu/_0368_ ) );
AOI221_X4 \myexu/_3328_ ( .A(\myexu/_0366_ ), .B1(\myexu/_0367_ ), .B2(\myexu/_2119_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0368_ ), .ZN(\myexu/_0369_ ) );
AND3_X1 \myexu/_3329_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1962_ ), .A3(\myexu/_2504_ ), .ZN(\myexu/_0370_ ) );
AOI221_X4 \myexu/_3330_ ( .A(\myexu/_0365_ ), .B1(\myexu/_1968_ ), .B2(\myexu/_0369_ ), .C1(\myexu/_2192_ ), .C2(\myexu/_0370_ ), .ZN(\myexu/_0371_ ) );
AOI21_X1 \myexu/_3331_ ( .A(\myexu/_2375_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_2046_ ), .ZN(\myexu/_0372_ ) );
NOR2_X1 \myexu/_3332_ ( .A1(\myexu/_0371_ ), .A2(\myexu/_0372_ ), .ZN(\myexu/_0099_ ) );
OAI21_X1 \myexu/_3333_ ( .A(\myexu/_2376_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_0373_ ) );
NAND4_X1 \myexu/_3334_ ( .A1(\myexu/_1979_ ), .A2(\myexu/_2001_ ), .A3(\myexu/_2473_ ), .A4(\myexu/_2003_ ), .ZN(\myexu/_0374_ ) );
OR2_X1 \myexu/_3335_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0309_ ), .ZN(\myexu/_0375_ ) );
OAI221_X1 \myexu/_3336_ ( .A(\myexu/_0375_ ), .B1(\myexu/_2441_ ), .B2(fanout_net_7 ), .C1(\myexu/_2114_ ), .C2(\myexu/_2505_ ), .ZN(\myexu/_0376_ ) );
NAND3_X1 \myexu/_3337_ ( .A1(\myexu/_2115_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2505_ ), .ZN(\myexu/_0377_ ) );
AOI21_X1 \myexu/_3338_ ( .A(\myexu/_2140_ ), .B1(\myexu/_0376_ ), .B2(\myexu/_0377_ ), .ZN(\myexu/_0378_ ) );
AOI21_X1 \myexu/_3339_ ( .A(\myexu/_0378_ ), .B1(\myexu/_2274_ ), .B2(\myexu/_2133_ ), .ZN(\myexu/_0379_ ) );
OAI211_X2 \myexu/_3340_ ( .A(\myexu/_0373_ ), .B(\myexu/_0374_ ), .C1(\myexu/_0379_ ), .C2(\myexu/_2072_ ), .ZN(\myexu/_0100_ ) );
AOI211_X4 \myexu/_3341_ ( .A(fanout_net_5 ), .B(\myexu/_1982_ ), .C1(\myexu/_2474_ ), .C2(\myexu/_1959_ ), .ZN(\myexu/_0380_ ) );
NAND3_X1 \myexu/_3342_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_2528_ ), .A3(\myexu/_2275_ ), .ZN(\myexu/_0381_ ) );
NAND2_X1 \myexu/_3343_ ( .A1(\myexu/_0380_ ), .A2(\myexu/_0381_ ), .ZN(\myexu/_0382_ ) );
NOR2_X1 \myexu/_3344_ ( .A1(\myexu/_2119_ ), .A2(\myexu/_0310_ ), .ZN(\myexu/_0383_ ) );
INV_X1 \myexu/_3345_ ( .A(\myexu/_2442_ ), .ZN(\myexu/_0384_ ) );
INV_X1 \myexu/_3346_ ( .A(\myexu/_2506_ ), .ZN(\myexu/_0385_ ) );
AOI221_X4 \myexu/_3347_ ( .A(\myexu/_0383_ ), .B1(\myexu/_0384_ ), .B2(\myexu/_2119_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0385_ ), .ZN(\myexu/_0386_ ) );
AND3_X1 \myexu/_3348_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1962_ ), .A3(\myexu/_2506_ ), .ZN(\myexu/_0387_ ) );
AOI221_X4 \myexu/_3349_ ( .A(\myexu/_0382_ ), .B1(\myexu/_1968_ ), .B2(\myexu/_0386_ ), .C1(\myexu/_2192_ ), .C2(\myexu/_0387_ ), .ZN(\myexu/_0388_ ) );
AOI21_X1 \myexu/_3350_ ( .A(\myexu/_2377_ ), .B1(\myexu/_2045_ ), .B2(\myexu/_2046_ ), .ZN(\myexu/_0389_ ) );
NOR2_X1 \myexu/_3351_ ( .A1(\myexu/_0388_ ), .A2(\myexu/_0389_ ), .ZN(\myexu/_0101_ ) );
AOI221_X4 \myexu/_3352_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2475_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2276_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_0390_ ) );
NOR2_X1 \myexu/_3353_ ( .A1(\myexu/_2120_ ), .A2(\myexu/_0311_ ), .ZN(\myexu/_0391_ ) );
INV_X1 \myexu/_3354_ ( .A(\myexu/_2443_ ), .ZN(\myexu/_0392_ ) );
INV_X1 \myexu/_3355_ ( .A(\myexu/_2507_ ), .ZN(\myexu/_0393_ ) );
AOI221_X4 \myexu/_3356_ ( .A(\myexu/_0391_ ), .B1(\myexu/_0392_ ), .B2(\myexu/_2127_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0393_ ), .ZN(\myexu/_0394_ ) );
NAND2_X1 \myexu/_3357_ ( .A1(\myexu/_0394_ ), .A2(\myexu/_2049_ ), .ZN(\myexu/_0395_ ) );
NAND3_X1 \myexu/_3358_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2507_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_0396_ ) );
NAND3_X1 \myexu/_3359_ ( .A1(\myexu/_0390_ ), .A2(\myexu/_0395_ ), .A3(\myexu/_0396_ ), .ZN(\myexu/_0397_ ) );
OR2_X1 \myexu/_3360_ ( .A1(\myexu/_1975_ ), .A2(\myexu/_2378_ ), .ZN(\myexu/_0398_ ) );
AND2_X1 \myexu/_3361_ ( .A1(\myexu/_0397_ ), .A2(\myexu/_0398_ ), .ZN(\myexu/_0102_ ) );
NOR2_X1 \myexu/_3362_ ( .A1(\myexu/_2119_ ), .A2(\myexu/_0312_ ), .ZN(\myexu/_0399_ ) );
INV_X1 \myexu/_3363_ ( .A(\myexu/_2444_ ), .ZN(\myexu/_0400_ ) );
INV_X1 \myexu/_3364_ ( .A(\myexu/_2508_ ), .ZN(\myexu/_0401_ ) );
AOI221_X4 \myexu/_3365_ ( .A(\myexu/_0399_ ), .B1(\myexu/_0400_ ), .B2(\myexu/_2120_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0401_ ), .ZN(\myexu/_0402_ ) );
AND3_X1 \myexu/_3366_ ( .A1(\myexu/_2113_ ), .A2(\myexu/_2524_ ), .A3(\myexu/_2508_ ), .ZN(\myexu/_0403_ ) );
OAI21_X1 \myexu/_3367_ ( .A(\myexu/_1968_ ), .B1(\myexu/_0402_ ), .B2(\myexu/_0403_ ), .ZN(\myexu/_0404_ ) );
INV_X1 \myexu/_3368_ ( .A(\myexu/_2476_ ), .ZN(\myexu/_0405_ ) );
INV_X1 \myexu/_3369_ ( .A(\myexu/_2277_ ), .ZN(\myexu/_0406_ ) );
OAI221_X1 \myexu/_3370_ ( .A(\myexu/_0404_ ), .B1(\myexu/_0405_ ), .B2(\myexu/_2057_ ), .C1(\myexu/_0406_ ), .C2(\myexu/_2030_ ), .ZN(\myexu/_0407_ ) );
MUX2_X1 \myexu/_3371_ ( .A(\myexu/_2379_ ), .B(\myexu/_0407_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0103_ ) );
AOI221_X4 \myexu/_3372_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2477_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2278_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_0408_ ) );
NOR2_X1 \myexu/_3373_ ( .A1(\myexu/_2120_ ), .A2(\myexu/_0313_ ), .ZN(\myexu/_0409_ ) );
INV_X1 \myexu/_3374_ ( .A(\myexu/_2445_ ), .ZN(\myexu/_0410_ ) );
INV_X1 \myexu/_3375_ ( .A(\myexu/_2509_ ), .ZN(\myexu/_0411_ ) );
AOI221_X4 \myexu/_3376_ ( .A(\myexu/_0409_ ), .B1(\myexu/_0410_ ), .B2(\myexu/_2127_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0411_ ), .ZN(\myexu/_0412_ ) );
NAND2_X1 \myexu/_3377_ ( .A1(\myexu/_0412_ ), .A2(\myexu/_2049_ ), .ZN(\myexu/_0413_ ) );
NAND3_X1 \myexu/_3378_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2509_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_0414_ ) );
NAND3_X1 \myexu/_3379_ ( .A1(\myexu/_0408_ ), .A2(\myexu/_0413_ ), .A3(\myexu/_0414_ ), .ZN(\myexu/_0415_ ) );
OR2_X1 \myexu/_3380_ ( .A1(\myexu/_1975_ ), .A2(\myexu/_2380_ ), .ZN(\myexu/_0416_ ) );
AND2_X1 \myexu/_3381_ ( .A1(\myexu/_0415_ ), .A2(\myexu/_0416_ ), .ZN(\myexu/_0104_ ) );
AOI21_X1 \myexu/_3382_ ( .A(\myexu/_2381_ ), .B1(\myexu/_1988_ ), .B2(\myexu/_2001_ ), .ZN(\myexu/_0417_ ) );
INV_X1 \myexu/_3383_ ( .A(\myexu/_2478_ ), .ZN(\myexu/_0418_ ) );
INV_X1 \myexu/_3384_ ( .A(\myexu/_2279_ ), .ZN(\myexu/_0419_ ) );
OAI221_X1 \myexu/_3385_ ( .A(\myexu/_2012_ ), .B1(\myexu/_0418_ ), .B2(\myexu/_2033_ ), .C1(\myexu/_2031_ ), .C2(\myexu/_0419_ ), .ZN(\myexu/_0420_ ) );
AND3_X1 \myexu/_3386_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2510_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_0421_ ) );
NOR2_X1 \myexu/_3387_ ( .A1(\myexu/_0420_ ), .A2(\myexu/_0421_ ), .ZN(\myexu/_0422_ ) );
INV_X1 \myexu/_3388_ ( .A(\myexu/_2446_ ), .ZN(\myexu/_0423_ ) );
NAND2_X1 \myexu/_3389_ ( .A1(\myexu/_0423_ ), .A2(\myexu/_2121_ ), .ZN(\myexu/_0424_ ) );
OAI221_X1 \myexu/_3390_ ( .A(\myexu/_0424_ ), .B1(\myexu/_0314_ ), .B2(\myexu/_2121_ ), .C1(\myexu/_2115_ ), .C2(\myexu/_2510_ ), .ZN(\myexu/_0425_ ) );
OR2_X1 \myexu/_3391_ ( .A1(\myexu/_0425_ ), .A2(\myexu/_2140_ ), .ZN(\myexu/_0426_ ) );
AOI21_X1 \myexu/_3392_ ( .A(\myexu/_0417_ ), .B1(\myexu/_0422_ ), .B2(\myexu/_0426_ ), .ZN(\myexu/_0105_ ) );
AOI21_X1 \myexu/_3393_ ( .A(\myexu/_2382_ ), .B1(\myexu/_1988_ ), .B2(\myexu/_2001_ ), .ZN(\myexu/_0427_ ) );
AOI211_X4 \myexu/_3394_ ( .A(fanout_net_5 ), .B(\myexu/_1982_ ), .C1(\myexu/_2479_ ), .C2(\myexu/_1961_ ), .ZN(\myexu/_0428_ ) );
NAND3_X1 \myexu/_3395_ ( .A1(\myexu/_2033_ ), .A2(\myexu/_2528_ ), .A3(\myexu/_2280_ ), .ZN(\myexu/_0429_ ) );
NAND2_X1 \myexu/_3396_ ( .A1(\myexu/_0428_ ), .A2(\myexu/_0429_ ), .ZN(\myexu/_0430_ ) );
INV_X1 \myexu/_3397_ ( .A(\myexu/_0315_ ), .ZN(\myexu/_0431_ ) );
NAND2_X1 \myexu/_3398_ ( .A1(\myexu/_0431_ ), .A2(fanout_net_7 ), .ZN(\myexu/_0432_ ) );
OAI221_X1 \myexu/_3399_ ( .A(\myexu/_0432_ ), .B1(\myexu/_2447_ ), .B2(fanout_net_7 ), .C1(\myexu/_2115_ ), .C2(\myexu/_2511_ ), .ZN(\myexu/_0433_ ) );
NOR2_X1 \myexu/_3400_ ( .A1(\myexu/_2140_ ), .A2(\myexu/_0433_ ), .ZN(\myexu/_0434_ ) );
NOR2_X1 \myexu/_3401_ ( .A1(\myexu/_0430_ ), .A2(\myexu/_0434_ ), .ZN(\myexu/_0435_ ) );
AND3_X1 \myexu/_3402_ ( .A1(\myexu/_2032_ ), .A2(\myexu/_1962_ ), .A3(\myexu/_2511_ ), .ZN(\myexu/_0436_ ) );
NAND2_X1 \myexu/_3403_ ( .A1(\myexu/_0436_ ), .A2(\myexu/_2109_ ), .ZN(\myexu/_0437_ ) );
AOI21_X1 \myexu/_3404_ ( .A(\myexu/_0427_ ), .B1(\myexu/_0435_ ), .B2(\myexu/_0437_ ), .ZN(\myexu/_0106_ ) );
AOI21_X1 \myexu/_3405_ ( .A(\myexu/_2383_ ), .B1(\myexu/_1988_ ), .B2(\myexu/_2001_ ), .ZN(\myexu/_0438_ ) );
INV_X1 \myexu/_3406_ ( .A(\myexu/_2480_ ), .ZN(\myexu/_0439_ ) );
BUF_X4 \myexu/_3407_ ( .A(\myexu/_2030_ ), .Z(\myexu/_0440_ ) );
INV_X1 \myexu/_3408_ ( .A(\myexu/_2281_ ), .ZN(\myexu/_0441_ ) );
OAI221_X1 \myexu/_3409_ ( .A(\myexu/_2082_ ), .B1(\myexu/_0439_ ), .B2(\myexu/_2033_ ), .C1(\myexu/_0440_ ), .C2(\myexu/_0441_ ), .ZN(\myexu/_0442_ ) );
NAND3_X1 \myexu/_3410_ ( .A1(\myexu/_2033_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2512_ ), .ZN(\myexu/_0443_ ) );
INV_X1 \myexu/_3411_ ( .A(\myexu/_2108_ ), .ZN(\myexu/_0444_ ) );
NOR2_X1 \myexu/_3412_ ( .A1(\myexu/_0443_ ), .A2(\myexu/_0444_ ), .ZN(\myexu/_0445_ ) );
NOR2_X1 \myexu/_3413_ ( .A1(\myexu/_0442_ ), .A2(\myexu/_0445_ ), .ZN(\myexu/_0446_ ) );
NOR2_X1 \myexu/_3414_ ( .A1(\myexu/_2153_ ), .A2(\myexu/_0316_ ), .ZN(\myexu/_0447_ ) );
INV_X1 \myexu/_3415_ ( .A(\myexu/_2448_ ), .ZN(\myexu/_0448_ ) );
INV_X1 \myexu/_3416_ ( .A(\myexu/_2512_ ), .ZN(\myexu/_0449_ ) );
AOI221_X4 \myexu/_3417_ ( .A(\myexu/_0447_ ), .B1(\myexu/_0448_ ), .B2(\myexu/_2121_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0449_ ), .ZN(\myexu/_0450_ ) );
NAND2_X1 \myexu/_3418_ ( .A1(\myexu/_0450_ ), .A2(\myexu/_1985_ ), .ZN(\myexu/_0451_ ) );
AOI21_X1 \myexu/_3419_ ( .A(\myexu/_0438_ ), .B1(\myexu/_0446_ ), .B2(\myexu/_0451_ ), .ZN(\myexu/_0107_ ) );
AOI21_X1 \myexu/_3420_ ( .A(\myexu/_2385_ ), .B1(\myexu/_1988_ ), .B2(\myexu/_2001_ ), .ZN(\myexu/_0452_ ) );
AOI211_X4 \myexu/_3421_ ( .A(fanout_net_5 ), .B(\myexu/_1982_ ), .C1(\myexu/_2482_ ), .C2(\myexu/_1961_ ), .ZN(\myexu/_0453_ ) );
NAND3_X1 \myexu/_3422_ ( .A1(\myexu/_2033_ ), .A2(\myexu/_2528_ ), .A3(\myexu/_2283_ ), .ZN(\myexu/_0454_ ) );
NAND2_X1 \myexu/_3423_ ( .A1(\myexu/_0453_ ), .A2(\myexu/_0454_ ), .ZN(\myexu/_0455_ ) );
INV_X1 \myexu/_3424_ ( .A(\myexu/_0318_ ), .ZN(\myexu/_0456_ ) );
NAND2_X1 \myexu/_3425_ ( .A1(\myexu/_0456_ ), .A2(fanout_net_7 ), .ZN(\myexu/_0457_ ) );
OAI221_X1 \myexu/_3426_ ( .A(\myexu/_0457_ ), .B1(\myexu/_2450_ ), .B2(fanout_net_7 ), .C1(\myexu/_2115_ ), .C2(\myexu/_2514_ ), .ZN(\myexu/_0458_ ) );
NOR2_X1 \myexu/_3427_ ( .A1(\myexu/_2140_ ), .A2(\myexu/_0458_ ), .ZN(\myexu/_0459_ ) );
NOR2_X1 \myexu/_3428_ ( .A1(\myexu/_0455_ ), .A2(\myexu/_0459_ ), .ZN(\myexu/_0460_ ) );
AND3_X1 \myexu/_3429_ ( .A1(\myexu/_2033_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2514_ ), .ZN(\myexu/_0461_ ) );
NAND2_X1 \myexu/_3430_ ( .A1(\myexu/_0461_ ), .A2(\myexu/_2109_ ), .ZN(\myexu/_0462_ ) );
AOI21_X1 \myexu/_3431_ ( .A(\myexu/_0452_ ), .B1(\myexu/_0460_ ), .B2(\myexu/_0462_ ), .ZN(\myexu/_0108_ ) );
AOI221_X4 \myexu/_3432_ ( .A(\myexu/_2071_ ), .B1(\myexu/_2483_ ), .B2(\myexu/_1960_ ), .C1(\myexu/_2284_ ), .C2(\myexu/_2070_ ), .ZN(\myexu/_0463_ ) );
NOR2_X1 \myexu/_3433_ ( .A1(\myexu/_2120_ ), .A2(\myexu/_0319_ ), .ZN(\myexu/_0464_ ) );
INV_X1 \myexu/_3434_ ( .A(\myexu/_2451_ ), .ZN(\myexu/_0465_ ) );
INV_X1 \myexu/_3435_ ( .A(\myexu/_2515_ ), .ZN(\myexu/_0466_ ) );
AOI221_X4 \myexu/_3436_ ( .A(\myexu/_0464_ ), .B1(\myexu/_0465_ ), .B2(\myexu/_2127_ ), .C1(\myexu/_2525_ ), .C2(\myexu/_0466_ ), .ZN(\myexu/_0467_ ) );
NAND2_X1 \myexu/_3437_ ( .A1(\myexu/_0467_ ), .A2(\myexu/_2049_ ), .ZN(\myexu/_0468_ ) );
NAND3_X1 \myexu/_3438_ ( .A1(\myexu/_2158_ ), .A2(\myexu/_2515_ ), .A3(\myexu/_2192_ ), .ZN(\myexu/_0469_ ) );
NAND3_X1 \myexu/_3439_ ( .A1(\myexu/_0463_ ), .A2(\myexu/_0468_ ), .A3(\myexu/_0469_ ), .ZN(\myexu/_0470_ ) );
OR2_X1 \myexu/_3440_ ( .A1(\myexu/_1975_ ), .A2(\myexu/_2386_ ), .ZN(\myexu/_0471_ ) );
AND2_X1 \myexu/_3441_ ( .A1(\myexu/_0470_ ), .A2(\myexu/_0471_ ), .ZN(\myexu/_0109_ ) );
INV_X1 \myexu/_3442_ ( .A(\myexu/_2065_ ), .ZN(\myexu/_0472_ ) );
AND2_X1 \myexu/_3443_ ( .A1(\myexu/_2085_ ), .A2(\myexu/_2100_ ), .ZN(\myexu/_0473_ ) );
INV_X1 \myexu/_3444_ ( .A(\myexu/_0473_ ), .ZN(\myexu/_0474_ ) );
NOR3_X1 \myexu/_3445_ ( .A1(\myexu/_0474_ ), .A2(\myexu/_2074_ ), .A3(\myexu/_2078_ ), .ZN(\myexu/_0475_ ) );
NAND2_X1 \myexu/_3446_ ( .A1(\myexu/_0472_ ), .A2(\myexu/_0475_ ), .ZN(\myexu/_0476_ ) );
NAND2_X1 \myexu/_3447_ ( .A1(\myexu/_2089_ ), .A2(\myexu/_0473_ ), .ZN(\myexu/_0477_ ) );
AND2_X1 \myexu/_3448_ ( .A1(\myexu/_2100_ ), .A2(\myexu/_2097_ ), .ZN(\myexu/_0478_ ) );
AOI21_X1 \myexu/_3449_ ( .A(\myexu/_0478_ ), .B1(\myexu/_2429_ ), .B2(\myexu/_0297_ ), .ZN(\myexu/_0479_ ) );
AND2_X1 \myexu/_3450_ ( .A1(\myexu/_0477_ ), .A2(\myexu/_0479_ ), .ZN(\myexu/_0480_ ) );
NAND2_X1 \myexu/_3451_ ( .A1(\myexu/_0476_ ), .A2(\myexu/_0480_ ), .ZN(\myexu/_0481_ ) );
XOR2_X1 \myexu/_3452_ ( .A(\myexu/_2430_ ), .B(\myexu/_0298_ ), .Z(\myexu/_0482_ ) );
XNOR2_X1 \myexu/_3453_ ( .A(\myexu/_0481_ ), .B(\myexu/_0482_ ), .ZN(\myexu/_0483_ ) );
NOR2_X1 \myexu/_3454_ ( .A1(\myexu/_0483_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0484_ ) );
MUX2_X1 \myexu/_3455_ ( .A(\myexu/_0258_ ), .B(\myexu/_0484_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0189_ ) );
NAND2_X1 \myexu/_3456_ ( .A1(\myexu/_0481_ ), .A2(\myexu/_0482_ ), .ZN(\myexu/_0485_ ) );
NAND2_X1 \myexu/_3457_ ( .A1(\myexu/_2430_ ), .A2(\myexu/_0298_ ), .ZN(\myexu/_0486_ ) );
AND2_X1 \myexu/_3458_ ( .A1(\myexu/_0485_ ), .A2(\myexu/_0486_ ), .ZN(\myexu/_0487_ ) );
AND2_X1 \myexu/_3459_ ( .A1(\myexu/_2431_ ), .A2(\myexu/_0299_ ), .ZN(\myexu/_0488_ ) );
NOR2_X1 \myexu/_3460_ ( .A1(\myexu/_2431_ ), .A2(\myexu/_0299_ ), .ZN(\myexu/_0489_ ) );
NOR2_X1 \myexu/_3461_ ( .A1(\myexu/_0488_ ), .A2(\myexu/_0489_ ), .ZN(\myexu/_0490_ ) );
XNOR2_X1 \myexu/_3462_ ( .A(\myexu/_0487_ ), .B(\myexu/_0490_ ), .ZN(\myexu/_0491_ ) );
AND2_X1 \myexu/_3463_ ( .A1(\myexu/_0491_ ), .A2(\myexu/_1979_ ), .ZN(\myexu/_0492_ ) );
MUX2_X1 \myexu/_3464_ ( .A(\myexu/_0259_ ), .B(\myexu/_0492_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0190_ ) );
AND2_X1 \myexu/_3465_ ( .A1(\myexu/_0482_ ), .A2(\myexu/_0490_ ), .ZN(\myexu/_0493_ ) );
AND2_X1 \myexu/_3466_ ( .A1(\myexu/_0481_ ), .A2(\myexu/_0493_ ), .ZN(\myexu/_0494_ ) );
INV_X1 \myexu/_3467_ ( .A(\myexu/_0488_ ), .ZN(\myexu/_0495_ ) );
AOI21_X1 \myexu/_3468_ ( .A(\myexu/_0489_ ), .B1(\myexu/_0495_ ), .B2(\myexu/_0486_ ), .ZN(\myexu/_0496_ ) );
XOR2_X1 \myexu/_3469_ ( .A(\myexu/_2432_ ), .B(\myexu/_0300_ ), .Z(\myexu/_0497_ ) );
OR3_X1 \myexu/_3470_ ( .A1(\myexu/_0494_ ), .A2(\myexu/_0496_ ), .A3(\myexu/_0497_ ), .ZN(\myexu/_0498_ ) );
OAI21_X1 \myexu/_3471_ ( .A(\myexu/_0497_ ), .B1(\myexu/_0494_ ), .B2(\myexu/_0496_ ), .ZN(\myexu/_0499_ ) );
AND3_X1 \myexu/_3472_ ( .A1(\myexu/_0498_ ), .A2(\myexu/_2207_ ), .A3(\myexu/_0499_ ), .ZN(\myexu/_0500_ ) );
MUX2_X1 \myexu/_3473_ ( .A(\myexu/_0260_ ), .B(\myexu/_0500_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0191_ ) );
AND2_X1 \myexu/_3474_ ( .A1(\myexu/_2432_ ), .A2(\myexu/_0300_ ), .ZN(\myexu/_0501_ ) );
INV_X1 \myexu/_3475_ ( .A(\myexu/_0501_ ), .ZN(\myexu/_0502_ ) );
NAND2_X1 \myexu/_3476_ ( .A1(\myexu/_0499_ ), .A2(\myexu/_0502_ ), .ZN(\myexu/_0503_ ) );
XOR2_X1 \myexu/_3477_ ( .A(\myexu/_2433_ ), .B(\myexu/_0301_ ), .Z(\myexu/_0504_ ) );
XNOR2_X1 \myexu/_3478_ ( .A(\myexu/_0503_ ), .B(\myexu/_0504_ ), .ZN(\myexu/_0505_ ) );
NOR2_X1 \myexu/_3479_ ( .A1(\myexu/_0505_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0506_ ) );
MUX2_X1 \myexu/_3480_ ( .A(\myexu/_0261_ ), .B(\myexu/_0506_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0192_ ) );
AND3_X1 \myexu/_3481_ ( .A1(\myexu/_0493_ ), .A2(\myexu/_0497_ ), .A3(\myexu/_0504_ ), .ZN(\myexu/_0507_ ) );
NAND3_X1 \myexu/_3482_ ( .A1(\myexu/_0472_ ), .A2(\myexu/_0475_ ), .A3(\myexu/_0507_ ), .ZN(\myexu/_0508_ ) );
NAND3_X1 \myexu/_3483_ ( .A1(\myexu/_0493_ ), .A2(\myexu/_0497_ ), .A3(\myexu/_0504_ ), .ZN(\myexu/_0509_ ) );
AOI21_X1 \myexu/_3484_ ( .A(\myexu/_0509_ ), .B1(\myexu/_0477_ ), .B2(\myexu/_0479_ ), .ZN(\myexu/_0510_ ) );
AND2_X1 \myexu/_3485_ ( .A1(\myexu/_2433_ ), .A2(\myexu/_0301_ ), .ZN(\myexu/_0511_ ) );
AND3_X1 \myexu/_3486_ ( .A1(\myexu/_0496_ ), .A2(\myexu/_0497_ ), .A3(\myexu/_0504_ ), .ZN(\myexu/_0512_ ) );
AND2_X1 \myexu/_3487_ ( .A1(\myexu/_0504_ ), .A2(\myexu/_0501_ ), .ZN(\myexu/_0513_ ) );
NOR4_X1 \myexu/_3488_ ( .A1(\myexu/_0510_ ), .A2(\myexu/_0511_ ), .A3(\myexu/_0512_ ), .A4(\myexu/_0513_ ), .ZN(\myexu/_0514_ ) );
AND2_X1 \myexu/_3489_ ( .A1(\myexu/_0508_ ), .A2(\myexu/_0514_ ), .ZN(\myexu/_0515_ ) );
XOR2_X1 \myexu/_3490_ ( .A(\myexu/_2434_ ), .B(\myexu/_0302_ ), .Z(\myexu/_0516_ ) );
XNOR2_X1 \myexu/_3491_ ( .A(\myexu/_0515_ ), .B(\myexu/_0516_ ), .ZN(\myexu/_0517_ ) );
AND2_X1 \myexu/_3492_ ( .A1(\myexu/_0517_ ), .A2(\myexu/_2207_ ), .ZN(\myexu/_0518_ ) );
MUX2_X1 \myexu/_3493_ ( .A(\myexu/_0262_ ), .B(\myexu/_0518_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0193_ ) );
NOR2_X1 \myexu/_3494_ ( .A1(\myexu/_2434_ ), .A2(\myexu/_0302_ ), .ZN(\myexu/_0519_ ) );
AND2_X1 \myexu/_3495_ ( .A1(\myexu/_2434_ ), .A2(\myexu/_0302_ ), .ZN(\myexu/_0520_ ) );
NOR3_X1 \myexu/_3496_ ( .A1(\myexu/_0515_ ), .A2(\myexu/_0519_ ), .A3(\myexu/_0520_ ), .ZN(\myexu/_0521_ ) );
OR2_X1 \myexu/_3497_ ( .A1(\myexu/_0521_ ), .A2(\myexu/_0520_ ), .ZN(\myexu/_0522_ ) );
AND2_X1 \myexu/_3498_ ( .A1(\myexu/_2435_ ), .A2(\myexu/_0303_ ), .ZN(\myexu/_0523_ ) );
NOR2_X1 \myexu/_3499_ ( .A1(\myexu/_2435_ ), .A2(\myexu/_0303_ ), .ZN(\myexu/_0524_ ) );
NOR2_X1 \myexu/_3500_ ( .A1(\myexu/_0523_ ), .A2(\myexu/_0524_ ), .ZN(\myexu/_0525_ ) );
XNOR2_X1 \myexu/_3501_ ( .A(\myexu/_0522_ ), .B(\myexu/_0525_ ), .ZN(\myexu/_0526_ ) );
NOR2_X1 \myexu/_3502_ ( .A1(\myexu/_0526_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0527_ ) );
MUX2_X1 \myexu/_3503_ ( .A(\myexu/_0263_ ), .B(\myexu/_0527_ ), .S(\myexu/_2205_ ), .Z(\myexu/_0194_ ) );
AND2_X1 \myexu/_3504_ ( .A1(\myexu/_0516_ ), .A2(\myexu/_0525_ ), .ZN(\myexu/_0528_ ) );
INV_X1 \myexu/_3505_ ( .A(\myexu/_0528_ ), .ZN(\myexu/_0529_ ) );
AOI21_X1 \myexu/_3506_ ( .A(\myexu/_0529_ ), .B1(\myexu/_0508_ ), .B2(\myexu/_0514_ ), .ZN(\myexu/_0530_ ) );
AOI21_X1 \myexu/_3507_ ( .A(\myexu/_0523_ ), .B1(\myexu/_0525_ ), .B2(\myexu/_0520_ ), .ZN(\myexu/_0531_ ) );
INV_X1 \myexu/_3508_ ( .A(\myexu/_0531_ ), .ZN(\myexu/_0532_ ) );
NOR2_X1 \myexu/_3509_ ( .A1(\myexu/_0530_ ), .A2(\myexu/_0532_ ), .ZN(\myexu/_0533_ ) );
XOR2_X1 \myexu/_3510_ ( .A(\myexu/_2436_ ), .B(\myexu/_0304_ ), .Z(\myexu/_0534_ ) );
XNOR2_X1 \myexu/_3511_ ( .A(\myexu/_0533_ ), .B(\myexu/_0534_ ), .ZN(\myexu/_0535_ ) );
AND2_X1 \myexu/_3512_ ( .A1(\myexu/_0535_ ), .A2(\myexu/_2207_ ), .ZN(\myexu/_0536_ ) );
BUF_X4 \myexu/_3513_ ( .A(\myexu/_1975_ ), .Z(\myexu/_0537_ ) );
MUX2_X1 \myexu/_3514_ ( .A(\myexu/_0264_ ), .B(\myexu/_0536_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0195_ ) );
OAI21_X1 \myexu/_3515_ ( .A(\myexu/_0534_ ), .B1(\myexu/_0530_ ), .B2(\myexu/_0532_ ), .ZN(\myexu/_0538_ ) );
NAND2_X1 \myexu/_3516_ ( .A1(\myexu/_2436_ ), .A2(\myexu/_0304_ ), .ZN(\myexu/_0539_ ) );
NAND2_X1 \myexu/_3517_ ( .A1(\myexu/_0538_ ), .A2(\myexu/_0539_ ), .ZN(\myexu/_0540_ ) );
XOR2_X1 \myexu/_3518_ ( .A(\myexu/_2437_ ), .B(\myexu/_0305_ ), .Z(\myexu/_0541_ ) );
XNOR2_X1 \myexu/_3519_ ( .A(\myexu/_0540_ ), .B(\myexu/_0541_ ), .ZN(\myexu/_0542_ ) );
NOR2_X1 \myexu/_3520_ ( .A1(\myexu/_0542_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0543_ ) );
MUX2_X1 \myexu/_3521_ ( .A(\myexu/_0265_ ), .B(\myexu/_0543_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0196_ ) );
AND2_X1 \myexu/_3522_ ( .A1(\myexu/_0534_ ), .A2(\myexu/_0541_ ), .ZN(\myexu/_0544_ ) );
AND2_X1 \myexu/_3523_ ( .A1(\myexu/_0544_ ), .A2(\myexu/_0528_ ), .ZN(\myexu/_0545_ ) );
INV_X1 \myexu/_3524_ ( .A(\myexu/_0545_ ), .ZN(\myexu/_0546_ ) );
AOI21_X1 \myexu/_3525_ ( .A(\myexu/_0546_ ), .B1(\myexu/_0508_ ), .B2(\myexu/_0514_ ), .ZN(\myexu/_0547_ ) );
INV_X1 \myexu/_3526_ ( .A(\myexu/_0547_ ), .ZN(\myexu/_0548_ ) );
AND2_X1 \myexu/_3527_ ( .A1(\myexu/_0532_ ), .A2(\myexu/_0544_ ), .ZN(\myexu/_0549_ ) );
AND2_X1 \myexu/_3528_ ( .A1(\myexu/_2437_ ), .A2(\myexu/_0305_ ), .ZN(\myexu/_0550_ ) );
AND3_X1 \myexu/_3529_ ( .A1(\myexu/_0541_ ), .A2(\myexu/_2436_ ), .A3(\myexu/_0304_ ), .ZN(\myexu/_0551_ ) );
NOR3_X1 \myexu/_3530_ ( .A1(\myexu/_0549_ ), .A2(\myexu/_0550_ ), .A3(\myexu/_0551_ ), .ZN(\myexu/_0552_ ) );
NAND2_X1 \myexu/_3531_ ( .A1(\myexu/_0548_ ), .A2(\myexu/_0552_ ), .ZN(\myexu/_0553_ ) );
XOR2_X1 \myexu/_3532_ ( .A(\myexu/_2439_ ), .B(\myexu/_0307_ ), .Z(\myexu/_0554_ ) );
XNOR2_X1 \myexu/_3533_ ( .A(\myexu/_0553_ ), .B(\myexu/_0554_ ), .ZN(\myexu/_0555_ ) );
NOR2_X1 \myexu/_3534_ ( .A1(\myexu/_0555_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0556_ ) );
MUX2_X1 \myexu/_3535_ ( .A(\myexu/_0267_ ), .B(\myexu/_0556_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0197_ ) );
AND2_X1 \myexu/_3536_ ( .A1(\myexu/_0553_ ), .A2(\myexu/_0554_ ), .ZN(\myexu/_0557_ ) );
AND2_X1 \myexu/_3537_ ( .A1(\myexu/_2439_ ), .A2(\myexu/_0307_ ), .ZN(\myexu/_0558_ ) );
OR2_X1 \myexu/_3538_ ( .A1(\myexu/_0557_ ), .A2(\myexu/_0558_ ), .ZN(\myexu/_0559_ ) );
XOR2_X1 \myexu/_3539_ ( .A(\myexu/_2440_ ), .B(\myexu/_0308_ ), .Z(\myexu/_0560_ ) );
XNOR2_X1 \myexu/_3540_ ( .A(\myexu/_0559_ ), .B(\myexu/_0560_ ), .ZN(\myexu/_0561_ ) );
NOR2_X1 \myexu/_3541_ ( .A1(\myexu/_0561_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0562_ ) );
MUX2_X1 \myexu/_3542_ ( .A(\myexu/_0268_ ), .B(\myexu/_0562_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0198_ ) );
AND2_X1 \myexu/_3543_ ( .A1(\myexu/_0554_ ), .A2(\myexu/_0560_ ), .ZN(\myexu/_0563_ ) );
NAND2_X1 \myexu/_3544_ ( .A1(\myexu/_0553_ ), .A2(\myexu/_0563_ ), .ZN(\myexu/_0564_ ) );
AND2_X1 \myexu/_3545_ ( .A1(\myexu/_0560_ ), .A2(\myexu/_0558_ ), .ZN(\myexu/_0565_ ) );
AOI21_X1 \myexu/_3546_ ( .A(\myexu/_0565_ ), .B1(\myexu/_2440_ ), .B2(\myexu/_0308_ ), .ZN(\myexu/_0566_ ) );
NAND2_X1 \myexu/_3547_ ( .A1(\myexu/_0564_ ), .A2(\myexu/_0566_ ), .ZN(\myexu/_0567_ ) );
XOR2_X1 \myexu/_3548_ ( .A(\myexu/_2441_ ), .B(\myexu/_0309_ ), .Z(\myexu/_0568_ ) );
XNOR2_X1 \myexu/_3549_ ( .A(\myexu/_0567_ ), .B(\myexu/_0568_ ), .ZN(\myexu/_0569_ ) );
NOR2_X1 \myexu/_3550_ ( .A1(\myexu/_0569_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0570_ ) );
MUX2_X1 \myexu/_3551_ ( .A(\myexu/_0269_ ), .B(\myexu/_0570_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0199_ ) );
AND2_X1 \myexu/_3552_ ( .A1(\myexu/_0567_ ), .A2(\myexu/_0568_ ), .ZN(\myexu/_0571_ ) );
AND2_X1 \myexu/_3553_ ( .A1(\myexu/_2441_ ), .A2(\myexu/_0309_ ), .ZN(\myexu/_0572_ ) );
OR2_X1 \myexu/_3554_ ( .A1(\myexu/_0571_ ), .A2(\myexu/_0572_ ), .ZN(\myexu/_0573_ ) );
XOR2_X1 \myexu/_3555_ ( .A(\myexu/_2442_ ), .B(\myexu/_0310_ ), .Z(\myexu/_0574_ ) );
XNOR2_X1 \myexu/_3556_ ( .A(\myexu/_0573_ ), .B(\myexu/_0574_ ), .ZN(\myexu/_0575_ ) );
NOR2_X1 \myexu/_3557_ ( .A1(\myexu/_0575_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0576_ ) );
MUX2_X1 \myexu/_3558_ ( .A(\myexu/_0270_ ), .B(\myexu/_0576_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0200_ ) );
AND2_X1 \myexu/_3559_ ( .A1(\myexu/_0568_ ), .A2(\myexu/_0574_ ), .ZN(\myexu/_0577_ ) );
AND2_X1 \myexu/_3560_ ( .A1(\myexu/_0563_ ), .A2(\myexu/_0577_ ), .ZN(\myexu/_0578_ ) );
NAND2_X1 \myexu/_3561_ ( .A1(\myexu/_0547_ ), .A2(\myexu/_0578_ ), .ZN(\myexu/_0579_ ) );
AND2_X1 \myexu/_3562_ ( .A1(\myexu/_0574_ ), .A2(\myexu/_0572_ ), .ZN(\myexu/_0580_ ) );
INV_X1 \myexu/_3563_ ( .A(\myexu/_0578_ ), .ZN(\myexu/_0581_ ) );
INV_X1 \myexu/_3564_ ( .A(\myexu/_0577_ ), .ZN(\myexu/_0582_ ) );
OAI22_X1 \myexu/_3565_ ( .A1(\myexu/_0552_ ), .A2(\myexu/_0581_ ), .B1(\myexu/_0566_ ), .B2(\myexu/_0582_ ), .ZN(\myexu/_0583_ ) );
AOI211_X4 \myexu/_3566_ ( .A(\myexu/_0580_ ), .B(\myexu/_0583_ ), .C1(\myexu/_2442_ ), .C2(\myexu/_0310_ ), .ZN(\myexu/_0584_ ) );
NAND2_X1 \myexu/_3567_ ( .A1(\myexu/_0579_ ), .A2(\myexu/_0584_ ), .ZN(\myexu/_0585_ ) );
XOR2_X1 \myexu/_3568_ ( .A(\myexu/_2443_ ), .B(\myexu/_0311_ ), .Z(\myexu/_0586_ ) );
INV_X1 \myexu/_3569_ ( .A(\myexu/_0586_ ), .ZN(\myexu/_0587_ ) );
XNOR2_X1 \myexu/_3570_ ( .A(\myexu/_0585_ ), .B(\myexu/_0587_ ), .ZN(\myexu/_0588_ ) );
AND2_X1 \myexu/_3571_ ( .A1(\myexu/_0588_ ), .A2(\myexu/_2207_ ), .ZN(\myexu/_0589_ ) );
MUX2_X1 \myexu/_3572_ ( .A(\myexu/_0271_ ), .B(\myexu/_0589_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0201_ ) );
AOI21_X1 \myexu/_3573_ ( .A(\myexu/_0587_ ), .B1(\myexu/_0579_ ), .B2(\myexu/_0584_ ), .ZN(\myexu/_0590_ ) );
AND2_X1 \myexu/_3574_ ( .A1(\myexu/_2443_ ), .A2(\myexu/_0311_ ), .ZN(\myexu/_0591_ ) );
OR2_X1 \myexu/_3575_ ( .A1(\myexu/_0590_ ), .A2(\myexu/_0591_ ), .ZN(\myexu/_0592_ ) );
XOR2_X1 \myexu/_3576_ ( .A(\myexu/_2444_ ), .B(\myexu/_0312_ ), .Z(\myexu/_0593_ ) );
XNOR2_X1 \myexu/_3577_ ( .A(\myexu/_0592_ ), .B(\myexu/_0593_ ), .ZN(\myexu/_0594_ ) );
NOR2_X1 \myexu/_3578_ ( .A1(\myexu/_0594_ ), .A2(\myexu/_2080_ ), .ZN(\myexu/_0595_ ) );
MUX2_X1 \myexu/_3579_ ( .A(\myexu/_0272_ ), .B(\myexu/_0595_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0202_ ) );
NAND3_X1 \myexu/_3580_ ( .A1(\myexu/_0585_ ), .A2(\myexu/_0586_ ), .A3(\myexu/_0593_ ), .ZN(\myexu/_0596_ ) );
AND2_X1 \myexu/_3581_ ( .A1(\myexu/_0593_ ), .A2(\myexu/_0591_ ), .ZN(\myexu/_0597_ ) );
AOI21_X1 \myexu/_3582_ ( .A(\myexu/_0597_ ), .B1(\myexu/_2444_ ), .B2(\myexu/_0312_ ), .ZN(\myexu/_0598_ ) );
NAND2_X1 \myexu/_3583_ ( .A1(\myexu/_0596_ ), .A2(\myexu/_0598_ ), .ZN(\myexu/_0599_ ) );
XOR2_X1 \myexu/_3584_ ( .A(\myexu/_2445_ ), .B(\myexu/_0313_ ), .Z(\myexu/_0600_ ) );
XNOR2_X1 \myexu/_3585_ ( .A(\myexu/_0599_ ), .B(\myexu/_0600_ ), .ZN(\myexu/_0601_ ) );
NOR2_X1 \myexu/_3586_ ( .A1(\myexu/_0601_ ), .A2(\myexu/_2033_ ), .ZN(\myexu/_0602_ ) );
MUX2_X1 \myexu/_3587_ ( .A(\myexu/_0273_ ), .B(\myexu/_0602_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0203_ ) );
AND2_X1 \myexu/_3588_ ( .A1(\myexu/_0599_ ), .A2(\myexu/_0600_ ), .ZN(\myexu/_0603_ ) );
AND2_X1 \myexu/_3589_ ( .A1(\myexu/_2445_ ), .A2(\myexu/_0313_ ), .ZN(\myexu/_0604_ ) );
OR2_X1 \myexu/_3590_ ( .A1(\myexu/_0603_ ), .A2(\myexu/_0604_ ), .ZN(\myexu/_0605_ ) );
XOR2_X1 \myexu/_3591_ ( .A(\myexu/_2446_ ), .B(\myexu/_0314_ ), .Z(\myexu/_0606_ ) );
XNOR2_X1 \myexu/_3592_ ( .A(\myexu/_0605_ ), .B(\myexu/_0606_ ), .ZN(\myexu/_0607_ ) );
NOR2_X1 \myexu/_3593_ ( .A1(\myexu/_0607_ ), .A2(\myexu/_2033_ ), .ZN(\myexu/_0608_ ) );
MUX2_X1 \myexu/_3594_ ( .A(\myexu/_0274_ ), .B(\myexu/_0608_ ), .S(\myexu/_0537_ ), .Z(\myexu/_0204_ ) );
NAND3_X1 \myexu/_3595_ ( .A1(\myexu/_0599_ ), .A2(\myexu/_0600_ ), .A3(\myexu/_0606_ ), .ZN(\myexu/_0609_ ) );
AND2_X1 \myexu/_3596_ ( .A1(\myexu/_0606_ ), .A2(\myexu/_0604_ ), .ZN(\myexu/_0610_ ) );
AOI21_X1 \myexu/_3597_ ( .A(\myexu/_0610_ ), .B1(\myexu/_2446_ ), .B2(\myexu/_0314_ ), .ZN(\myexu/_0611_ ) );
NAND2_X1 \myexu/_3598_ ( .A1(\myexu/_0609_ ), .A2(\myexu/_0611_ ), .ZN(\myexu/_0612_ ) );
XOR2_X1 \myexu/_3599_ ( .A(\myexu/_2447_ ), .B(\myexu/_0315_ ), .Z(\myexu/_0613_ ) );
XOR2_X1 \myexu/_3600_ ( .A(\myexu/_0612_ ), .B(\myexu/_0613_ ), .Z(\myexu/_0614_ ) );
AND2_X1 \myexu/_3601_ ( .A1(\myexu/_0614_ ), .A2(\myexu/_2207_ ), .ZN(\myexu/_0615_ ) );
BUF_X4 \myexu/_3602_ ( .A(\myexu/_1975_ ), .Z(\myexu/_0616_ ) );
MUX2_X1 \myexu/_3603_ ( .A(\myexu/_0275_ ), .B(\myexu/_0615_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0205_ ) );
NAND2_X1 \myexu/_3604_ ( .A1(\myexu/_0612_ ), .A2(\myexu/_0613_ ), .ZN(\myexu/_0617_ ) );
NAND2_X1 \myexu/_3605_ ( .A1(\myexu/_2447_ ), .A2(\myexu/_0315_ ), .ZN(\myexu/_0618_ ) );
NAND2_X1 \myexu/_3606_ ( .A1(\myexu/_0617_ ), .A2(\myexu/_0618_ ), .ZN(\myexu/_0619_ ) );
XNOR2_X1 \myexu/_3607_ ( .A(\myexu/_2448_ ), .B(\myexu/_0316_ ), .ZN(\myexu/_0620_ ) );
XNOR2_X1 \myexu/_3608_ ( .A(\myexu/_0619_ ), .B(\myexu/_0620_ ), .ZN(\myexu/_0621_ ) );
AND2_X1 \myexu/_3609_ ( .A1(\myexu/_0621_ ), .A2(\myexu/_2207_ ), .ZN(\myexu/_0622_ ) );
MUX2_X1 \myexu/_3610_ ( .A(\myexu/_0276_ ), .B(\myexu/_0622_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0206_ ) );
OAI21_X1 \myexu/_3611_ ( .A(\myexu/_0619_ ), .B1(\myexu/_2448_ ), .B2(\myexu/_0316_ ), .ZN(\myexu/_0623_ ) );
NAND2_X1 \myexu/_3612_ ( .A1(\myexu/_2448_ ), .A2(\myexu/_0316_ ), .ZN(\myexu/_0624_ ) );
NAND2_X1 \myexu/_3613_ ( .A1(\myexu/_0623_ ), .A2(\myexu/_0624_ ), .ZN(\myexu/_0625_ ) );
XOR2_X1 \myexu/_3614_ ( .A(\myexu/_2450_ ), .B(\myexu/_0318_ ), .Z(\myexu/_0626_ ) );
XOR2_X1 \myexu/_3615_ ( .A(\myexu/_0625_ ), .B(\myexu/_0626_ ), .Z(\myexu/_0627_ ) );
AND2_X1 \myexu/_3616_ ( .A1(\myexu/_0627_ ), .A2(\myexu/_2207_ ), .ZN(\myexu/_0628_ ) );
MUX2_X1 \myexu/_3617_ ( .A(\myexu/_0278_ ), .B(\myexu/_0628_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0207_ ) );
NAND2_X1 \myexu/_3618_ ( .A1(\myexu/_0625_ ), .A2(\myexu/_0626_ ), .ZN(\myexu/_0629_ ) );
NAND2_X1 \myexu/_3619_ ( .A1(\myexu/_2450_ ), .A2(\myexu/_0318_ ), .ZN(\myexu/_0630_ ) );
NAND2_X1 \myexu/_3620_ ( .A1(\myexu/_0629_ ), .A2(\myexu/_0630_ ), .ZN(\myexu/_0631_ ) );
XOR2_X1 \myexu/_3621_ ( .A(\myexu/_0319_ ), .B(\myexu/_2451_ ), .Z(\myexu/_0632_ ) );
XNOR2_X1 \myexu/_3622_ ( .A(\myexu/_0631_ ), .B(\myexu/_0632_ ), .ZN(\myexu/_0633_ ) );
NOR2_X1 \myexu/_3623_ ( .A1(\myexu/_0633_ ), .A2(\myexu/_2033_ ), .ZN(\myexu/_0634_ ) );
MUX2_X1 \myexu/_3624_ ( .A(\myexu/_0279_ ), .B(\myexu/_0634_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0208_ ) );
INV_X1 \myexu/_3625_ ( .A(\myexu/_2110_ ), .ZN(\myexu/_0635_ ) );
NOR2_X1 \myexu/_3626_ ( .A1(\myexu/_1962_ ), .A2(\myexu/_2529_ ), .ZN(\myexu/_0636_ ) );
INV_X1 \myexu/_3627_ ( .A(\myexu/_2530_ ), .ZN(\myexu/_0637_ ) );
AND2_X1 \myexu/_3628_ ( .A1(\myexu/_0636_ ), .A2(\myexu/_0637_ ), .ZN(\myexu/_0638_ ) );
INV_X2 \myexu/_3629_ ( .A(\myexu/_0638_ ), .ZN(\myexu/_0639_ ) );
BUF_X4 \myexu/_3630_ ( .A(\myexu/_0639_ ), .Z(\myexu/_0640_ ) );
AND2_X1 \myexu/_3631_ ( .A1(\myexu/_0023_ ), .A2(\myexu/_0448_ ), .ZN(\myexu/_0641_ ) );
INV_X1 \myexu/_3632_ ( .A(\myexu/_2447_ ), .ZN(\myexu/_0642_ ) );
AND2_X1 \myexu/_3633_ ( .A1(\myexu/_0022_ ), .A2(\myexu/_0642_ ), .ZN(\myexu/_0643_ ) );
NOR2_X1 \myexu/_3634_ ( .A1(\myexu/_0022_ ), .A2(\myexu/_0642_ ), .ZN(\myexu/_0644_ ) );
NOR2_X1 \myexu/_3635_ ( .A1(\myexu/_0023_ ), .A2(\myexu/_0448_ ), .ZN(\myexu/_0645_ ) );
NOR4_X1 \myexu/_3636_ ( .A1(\myexu/_0641_ ), .A2(\myexu/_0643_ ), .A3(\myexu/_0644_ ), .A4(\myexu/_0645_ ), .ZN(\myexu/_0646_ ) );
XNOR2_X1 \myexu/_3637_ ( .A(\myexu/_0003_ ), .B(\myexu/_2428_ ), .ZN(\myexu/_0647_ ) );
XNOR2_X1 \myexu/_3638_ ( .A(\myexu/_0004_ ), .B(\myexu/_2429_ ), .ZN(\myexu/_0648_ ) );
AND2_X1 \myexu/_3639_ ( .A1(\myexu/_0647_ ), .A2(\myexu/_0648_ ), .ZN(\myexu/_0649_ ) );
XNOR2_X1 \myexu/_3640_ ( .A(\myexu/_0033_ ), .B(\myexu/_2458_ ), .ZN(\myexu/_0650_ ) );
XNOR2_X1 \myexu/_3641_ ( .A(\myexu/_0032_ ), .B(\myexu/_2457_ ), .ZN(\myexu/_0651_ ) );
AND3_X1 \myexu/_3642_ ( .A1(\myexu/_0649_ ), .A2(\myexu/_0650_ ), .A3(\myexu/_0651_ ), .ZN(\myexu/_0652_ ) );
XNOR2_X1 \myexu/_3643_ ( .A(\myexu/_0008_ ), .B(\myexu/_2433_ ), .ZN(\myexu/_0653_ ) );
INV_X1 \myexu/_3644_ ( .A(\myexu/_0653_ ), .ZN(\myexu/_0654_ ) );
INV_X1 \myexu/_3645_ ( .A(\myexu/_2432_ ), .ZN(\myexu/_0655_ ) );
AND2_X1 \myexu/_3646_ ( .A1(\myexu/_0007_ ), .A2(\myexu/_0655_ ), .ZN(\myexu/_0656_ ) );
NOR2_X1 \myexu/_3647_ ( .A1(\myexu/_0007_ ), .A2(\myexu/_0655_ ), .ZN(\myexu/_0657_ ) );
NOR3_X1 \myexu/_3648_ ( .A1(\myexu/_0654_ ), .A2(\myexu/_0656_ ), .A3(\myexu/_0657_ ), .ZN(\myexu/_0658_ ) );
INV_X1 \myexu/_3649_ ( .A(\myexu/_2431_ ), .ZN(\myexu/_0659_ ) );
XNOR2_X1 \myexu/_3650_ ( .A(\myexu/_0006_ ), .B(\myexu/_0659_ ), .ZN(\myexu/_0660_ ) );
XNOR2_X1 \myexu/_3651_ ( .A(\myexu/_0005_ ), .B(\myexu/_2226_ ), .ZN(\myexu/_0661_ ) );
NOR2_X1 \myexu/_3652_ ( .A1(\myexu/_0660_ ), .A2(\myexu/_0661_ ), .ZN(\myexu/_0662_ ) );
AND3_X1 \myexu/_3653_ ( .A1(\myexu/_0652_ ), .A2(\myexu/_0658_ ), .A3(\myexu/_0662_ ), .ZN(\myexu/_0663_ ) );
INV_X1 \myexu/_3654_ ( .A(\myexu/_2427_ ), .ZN(\myexu/_0664_ ) );
NAND3_X1 \myexu/_3655_ ( .A1(\myexu/_1927_ ), .A2(\myexu/_2438_ ), .A3(\myexu/_1928_ ), .ZN(\myexu/_0665_ ) );
AND3_X1 \myexu/_3656_ ( .A1(\myexu/_0002_ ), .A2(\myexu/_0664_ ), .A3(\myexu/_0665_ ), .ZN(\myexu/_0666_ ) );
AOI21_X1 \myexu/_3657_ ( .A(\myexu/_2438_ ), .B1(\myexu/_1927_ ), .B2(\myexu/_1928_ ), .ZN(\myexu/_0667_ ) );
INV_X1 \myexu/_3658_ ( .A(\myexu/_2452_ ), .ZN(\myexu/_0668_ ) );
NOR2_X1 \myexu/_3659_ ( .A1(\myexu/_0027_ ), .A2(\myexu/_0668_ ), .ZN(\myexu/_0669_ ) );
NOR2_X1 \myexu/_3660_ ( .A1(\myexu/_0024_ ), .A2(\myexu/_2137_ ), .ZN(\myexu/_0670_ ) );
AND3_X1 \myexu/_3661_ ( .A1(\myexu/_1930_ ), .A2(\myexu/_1932_ ), .A3(\myexu/_0668_ ), .ZN(\myexu/_0671_ ) );
OR4_X2 \myexu/_3662_ ( .A1(\myexu/_0667_ ), .A2(\myexu/_0669_ ), .A3(\myexu/_0670_ ), .A4(\myexu/_0671_ ), .ZN(\myexu/_0672_ ) );
AOI211_X2 \myexu/_3663_ ( .A(\myexu/_0666_ ), .B(\myexu/_0672_ ), .C1(\myexu/_2137_ ), .C2(\myexu/_0024_ ), .ZN(\myexu/_0673_ ) );
NOR4_X1 \myexu/_3664_ ( .A1(\myexu/_0669_ ), .A2(\myexu/_2137_ ), .A3(\myexu/_0024_ ), .A4(\myexu/_0671_ ), .ZN(\myexu/_0674_ ) );
NOR3_X1 \myexu/_3665_ ( .A1(\myexu/_0673_ ), .A2(\myexu/_0669_ ), .A3(\myexu/_0674_ ), .ZN(\myexu/_0675_ ) );
XNOR2_X1 \myexu/_3666_ ( .A(\myexu/_0030_ ), .B(\myexu/_2455_ ), .ZN(\myexu/_0676_ ) );
XNOR2_X1 \myexu/_3667_ ( .A(\myexu/_0029_ ), .B(\myexu/_2454_ ), .ZN(\myexu/_0677_ ) );
XNOR2_X1 \myexu/_3668_ ( .A(\myexu/_0028_ ), .B(\myexu/_2453_ ), .ZN(\myexu/_0678_ ) );
XNOR2_X1 \myexu/_3669_ ( .A(\myexu/_0031_ ), .B(\myexu/_2456_ ), .ZN(\myexu/_0679_ ) );
NAND4_X1 \myexu/_3670_ ( .A1(\myexu/_0676_ ), .A2(\myexu/_0677_ ), .A3(\myexu/_0678_ ), .A4(\myexu/_0679_ ), .ZN(\myexu/_0680_ ) );
NOR2_X1 \myexu/_3671_ ( .A1(\myexu/_0675_ ), .A2(\myexu/_0680_ ), .ZN(\myexu/_0681_ ) );
INV_X1 \myexu/_3672_ ( .A(\myexu/_2453_ ), .ZN(\myexu/_0682_ ) );
INV_X1 \myexu/_3673_ ( .A(\myexu/_2454_ ), .ZN(\myexu/_0683_ ) );
AOI211_X4 \myexu/_3674_ ( .A(\myexu/_0682_ ), .B(\myexu/_0028_ ), .C1(\myexu/_0683_ ), .C2(\myexu/_0029_ ), .ZN(\myexu/_0684_ ) );
NOR2_X1 \myexu/_3675_ ( .A1(\myexu/_0029_ ), .A2(\myexu/_0683_ ), .ZN(\myexu/_0685_ ) );
OAI211_X2 \myexu/_3676_ ( .A(\myexu/_0679_ ), .B(\myexu/_0676_ ), .C1(\myexu/_0684_ ), .C2(\myexu/_0685_ ), .ZN(\myexu/_0686_ ) );
NOR2_X1 \myexu/_3677_ ( .A1(\myexu/_0030_ ), .A2(\myexu/_2171_ ), .ZN(\myexu/_0687_ ) );
NAND2_X1 \myexu/_3678_ ( .A1(\myexu/_0679_ ), .A2(\myexu/_0687_ ), .ZN(\myexu/_0688_ ) );
OAI211_X2 \myexu/_3679_ ( .A(\myexu/_0686_ ), .B(\myexu/_0688_ ), .C1(\myexu/_2181_ ), .C2(\myexu/_0031_ ), .ZN(\myexu/_0689_ ) );
OAI21_X1 \myexu/_3680_ ( .A(\myexu/_0663_ ), .B1(\myexu/_0681_ ), .B2(\myexu/_0689_ ), .ZN(\myexu/_0690_ ) );
NOR3_X1 \myexu/_3681_ ( .A1(\myexu/_0660_ ), .A2(\myexu/_2226_ ), .A3(\myexu/_0005_ ), .ZN(\myexu/_0691_ ) );
NOR2_X1 \myexu/_3682_ ( .A1(\myexu/_0006_ ), .A2(\myexu/_0659_ ), .ZN(\myexu/_0692_ ) );
OAI21_X1 \myexu/_3683_ ( .A(\myexu/_0658_ ), .B1(\myexu/_0691_ ), .B2(\myexu/_0692_ ), .ZN(\myexu/_0693_ ) );
AND3_X1 \myexu/_3684_ ( .A1(\myexu/_1937_ ), .A2(\myexu/_2433_ ), .A3(\myexu/_1938_ ), .ZN(\myexu/_0694_ ) );
AOI21_X1 \myexu/_3685_ ( .A(\myexu/_0694_ ), .B1(\myexu/_0653_ ), .B2(\myexu/_0657_ ), .ZN(\myexu/_0695_ ) );
NOR2_X1 \myexu/_3686_ ( .A1(\myexu/_0033_ ), .A2(\myexu/_2197_ ), .ZN(\myexu/_0696_ ) );
INV_X1 \myexu/_3687_ ( .A(\myexu/_2457_ ), .ZN(\myexu/_0697_ ) );
AOI211_X4 \myexu/_3688_ ( .A(\myexu/_0697_ ), .B(\myexu/_0032_ ), .C1(\myexu/_2197_ ), .C2(\myexu/_0033_ ), .ZN(\myexu/_0698_ ) );
OAI21_X1 \myexu/_3689_ ( .A(\myexu/_0649_ ), .B1(\myexu/_0696_ ), .B2(\myexu/_0698_ ), .ZN(\myexu/_0699_ ) );
INV_X1 \myexu/_3690_ ( .A(\myexu/_2429_ ), .ZN(\myexu/_0700_ ) );
NOR2_X1 \myexu/_3691_ ( .A1(\myexu/_0004_ ), .A2(\myexu/_0700_ ), .ZN(\myexu/_0701_ ) );
NOR2_X1 \myexu/_3692_ ( .A1(\myexu/_0003_ ), .A2(\myexu/_2210_ ), .ZN(\myexu/_0702_ ) );
AOI21_X1 \myexu/_3693_ ( .A(\myexu/_0701_ ), .B1(\myexu/_0648_ ), .B2(\myexu/_0702_ ), .ZN(\myexu/_0703_ ) );
NAND2_X1 \myexu/_3694_ ( .A1(\myexu/_0699_ ), .A2(\myexu/_0703_ ), .ZN(\myexu/_0704_ ) );
NAND3_X1 \myexu/_3695_ ( .A1(\myexu/_0704_ ), .A2(\myexu/_0658_ ), .A3(\myexu/_0662_ ), .ZN(\myexu/_0705_ ) );
NAND4_X1 \myexu/_3696_ ( .A1(\myexu/_0690_ ), .A2(\myexu/_0693_ ), .A3(\myexu/_0695_ ), .A4(\myexu/_0705_ ), .ZN(\myexu/_0706_ ) );
XNOR2_X1 \myexu/_3697_ ( .A(\myexu/_0011_ ), .B(\myexu/_0342_ ), .ZN(\myexu/_0707_ ) );
AND2_X1 \myexu/_3698_ ( .A1(\myexu/_0012_ ), .A2(\myexu/_0348_ ), .ZN(\myexu/_0708_ ) );
NOR2_X1 \myexu/_3699_ ( .A1(\myexu/_0012_ ), .A2(\myexu/_0348_ ), .ZN(\myexu/_0709_ ) );
NOR3_X1 \myexu/_3700_ ( .A1(\myexu/_0707_ ), .A2(\myexu/_0708_ ), .A3(\myexu/_0709_ ), .ZN(\myexu/_0710_ ) );
XNOR2_X1 \myexu/_3701_ ( .A(\myexu/_0016_ ), .B(\myexu/_2441_ ), .ZN(\myexu/_0711_ ) );
XNOR2_X1 \myexu/_3702_ ( .A(\myexu/_0017_ ), .B(\myexu/_2442_ ), .ZN(\myexu/_0712_ ) );
AND2_X1 \myexu/_3703_ ( .A1(\myexu/_0711_ ), .A2(\myexu/_0712_ ), .ZN(\myexu/_0713_ ) );
INV_X1 \myexu/_3704_ ( .A(\myexu/_2439_ ), .ZN(\myexu/_0714_ ) );
XNOR2_X1 \myexu/_3705_ ( .A(\myexu/_0014_ ), .B(\myexu/_0714_ ), .ZN(\myexu/_0715_ ) );
NOR2_X1 \myexu/_3706_ ( .A1(\myexu/_0015_ ), .A2(\myexu/_0367_ ), .ZN(\myexu/_0716_ ) );
AND2_X1 \myexu/_3707_ ( .A1(\myexu/_0015_ ), .A2(\myexu/_0367_ ), .ZN(\myexu/_0717_ ) );
NOR3_X1 \myexu/_3708_ ( .A1(\myexu/_0715_ ), .A2(\myexu/_0716_ ), .A3(\myexu/_0717_ ), .ZN(\myexu/_0718_ ) );
OR3_X1 \myexu/_3709_ ( .A1(\myexu/_1940_ ), .A2(\myexu/_2434_ ), .A3(\myexu/_1941_ ), .ZN(\myexu/_0719_ ) );
NAND4_X1 \myexu/_3710_ ( .A1(\myexu/_0710_ ), .A2(\myexu/_0713_ ), .A3(\myexu/_0718_ ), .A4(\myexu/_0719_ ), .ZN(\myexu/_0720_ ) );
AOI21_X1 \myexu/_3711_ ( .A(\myexu/_2435_ ), .B1(\myexu/_1942_ ), .B2(\myexu/_1943_ ), .ZN(\myexu/_0721_ ) );
NOR2_X1 \myexu/_3712_ ( .A1(\myexu/_0010_ ), .A2(\myexu/_0333_ ), .ZN(\myexu/_0722_ ) );
INV_X1 \myexu/_3713_ ( .A(\myexu/_2434_ ), .ZN(\myexu/_0723_ ) );
NOR2_X1 \myexu/_3714_ ( .A1(\myexu/_0009_ ), .A2(\myexu/_0723_ ), .ZN(\myexu/_0724_ ) );
NOR4_X1 \myexu/_3715_ ( .A1(\myexu/_0720_ ), .A2(\myexu/_0721_ ), .A3(\myexu/_0722_ ), .A4(\myexu/_0724_ ), .ZN(\myexu/_0725_ ) );
NAND2_X1 \myexu/_3716_ ( .A1(\myexu/_0706_ ), .A2(\myexu/_0725_ ), .ZN(\myexu/_0726_ ) );
INV_X1 \myexu/_3717_ ( .A(\myexu/_2441_ ), .ZN(\myexu/_0727_ ) );
AOI211_X4 \myexu/_3718_ ( .A(\myexu/_0727_ ), .B(\myexu/_0016_ ), .C1(\myexu/_0384_ ), .C2(\myexu/_0017_ ), .ZN(\myexu/_0728_ ) );
NOR2_X1 \myexu/_3719_ ( .A1(\myexu/_0017_ ), .A2(\myexu/_0384_ ), .ZN(\myexu/_0729_ ) );
NOR2_X1 \myexu/_3720_ ( .A1(\myexu/_0728_ ), .A2(\myexu/_0729_ ), .ZN(\myexu/_0730_ ) );
NOR4_X1 \myexu/_3721_ ( .A1(\myexu/_0717_ ), .A2(\myexu/_0716_ ), .A3(\myexu/_0714_ ), .A4(\myexu/_0014_ ), .ZN(\myexu/_0731_ ) );
OAI21_X1 \myexu/_3722_ ( .A(\myexu/_0713_ ), .B1(\myexu/_0731_ ), .B2(\myexu/_0716_ ), .ZN(\myexu/_0732_ ) );
AND3_X1 \myexu/_3723_ ( .A1(\myexu/_0718_ ), .A2(\myexu/_0712_ ), .A3(\myexu/_0711_ ), .ZN(\myexu/_0733_ ) );
NOR4_X1 \myexu/_3724_ ( .A1(\myexu/_0722_ ), .A2(\myexu/_0721_ ), .A3(\myexu/_0009_ ), .A4(\myexu/_0723_ ), .ZN(\myexu/_0734_ ) );
OAI21_X1 \myexu/_3725_ ( .A(\myexu/_0710_ ), .B1(\myexu/_0722_ ), .B2(\myexu/_0734_ ), .ZN(\myexu/_0735_ ) );
OAI21_X1 \myexu/_3726_ ( .A(\myexu/_0735_ ), .B1(\myexu/_0348_ ), .B2(\myexu/_0012_ ), .ZN(\myexu/_0736_ ) );
NOR3_X1 \myexu/_3727_ ( .A1(\myexu/_0708_ ), .A2(\myexu/_0342_ ), .A3(\myexu/_0011_ ), .ZN(\myexu/_0737_ ) );
OAI21_X1 \myexu/_3728_ ( .A(\myexu/_0733_ ), .B1(\myexu/_0736_ ), .B2(\myexu/_0737_ ), .ZN(\myexu/_0738_ ) );
NAND4_X1 \myexu/_3729_ ( .A1(\myexu/_0726_ ), .A2(\myexu/_0730_ ), .A3(\myexu/_0732_ ), .A4(\myexu/_0738_ ), .ZN(\myexu/_0739_ ) );
XNOR2_X1 \myexu/_3730_ ( .A(\myexu/_0021_ ), .B(\myexu/_0423_ ), .ZN(\myexu/_0740_ ) );
AND2_X1 \myexu/_3731_ ( .A1(\myexu/_0020_ ), .A2(\myexu/_0410_ ), .ZN(\myexu/_0741_ ) );
NOR2_X1 \myexu/_3732_ ( .A1(\myexu/_0020_ ), .A2(\myexu/_0410_ ), .ZN(\myexu/_0742_ ) );
NOR3_X1 \myexu/_3733_ ( .A1(\myexu/_0740_ ), .A2(\myexu/_0741_ ), .A3(\myexu/_0742_ ), .ZN(\myexu/_0743_ ) );
XNOR2_X1 \myexu/_3734_ ( .A(\myexu/_0019_ ), .B(\myexu/_2444_ ), .ZN(\myexu/_0744_ ) );
XNOR2_X1 \myexu/_3735_ ( .A(\myexu/_0018_ ), .B(\myexu/_2443_ ), .ZN(\myexu/_0745_ ) );
AND4_X2 \myexu/_3736_ ( .A1(\myexu/_0739_ ), .A2(\myexu/_0743_ ), .A3(\myexu/_0744_ ), .A4(\myexu/_0745_ ), .ZN(\myexu/_0746_ ) );
OR2_X1 \myexu/_3737_ ( .A1(\myexu/_0018_ ), .A2(\myexu/_0392_ ), .ZN(\myexu/_0747_ ) );
AND2_X1 \myexu/_3738_ ( .A1(\myexu/_0019_ ), .A2(\myexu/_0400_ ), .ZN(\myexu/_0748_ ) );
NOR2_X1 \myexu/_3739_ ( .A1(\myexu/_0019_ ), .A2(\myexu/_0400_ ), .ZN(\myexu/_0749_ ) );
NOR3_X1 \myexu/_3740_ ( .A1(\myexu/_0747_ ), .A2(\myexu/_0748_ ), .A3(\myexu/_0749_ ), .ZN(\myexu/_0750_ ) );
OAI21_X1 \myexu/_3741_ ( .A(\myexu/_0743_ ), .B1(\myexu/_0750_ ), .B2(\myexu/_0749_ ), .ZN(\myexu/_0751_ ) );
OR3_X1 \myexu/_3742_ ( .A1(\myexu/_0740_ ), .A2(\myexu/_0410_ ), .A3(\myexu/_0020_ ), .ZN(\myexu/_0752_ ) );
OAI211_X2 \myexu/_3743_ ( .A(\myexu/_0751_ ), .B(\myexu/_0752_ ), .C1(\myexu/_0423_ ), .C2(\myexu/_0021_ ), .ZN(\myexu/_0753_ ) );
OAI21_X2 \myexu/_3744_ ( .A(\myexu/_0646_ ), .B1(\myexu/_0746_ ), .B2(\myexu/_0753_ ), .ZN(\myexu/_0754_ ) );
INV_X1 \myexu/_3745_ ( .A(\myexu/_2450_ ), .ZN(\myexu/_0755_ ) );
NOR2_X1 \myexu/_3746_ ( .A1(\myexu/_0644_ ), .A2(\myexu/_0645_ ), .ZN(\myexu/_0756_ ) );
OAI221_X2 \myexu/_3747_ ( .A(\myexu/_0754_ ), .B1(\myexu/_0755_ ), .B2(\myexu/_0025_ ), .C1(\myexu/_0641_ ), .C2(\myexu/_0756_ ), .ZN(\myexu/_0757_ ) );
NAND2_X1 \myexu/_3748_ ( .A1(\myexu/_0025_ ), .A2(\myexu/_0755_ ), .ZN(\myexu/_0758_ ) );
OAI211_X2 \myexu/_3749_ ( .A(\myexu/_0757_ ), .B(\myexu/_0758_ ), .C1(\myexu/_0465_ ), .C2(\myexu/_0026_ ), .ZN(\myexu/_0759_ ) );
NAND2_X1 \myexu/_3750_ ( .A1(\myexu/_0026_ ), .A2(\myexu/_0465_ ), .ZN(\myexu/_0760_ ) );
NAND2_X2 \myexu/_3751_ ( .A1(\myexu/_0759_ ), .A2(\myexu/_0760_ ), .ZN(\myexu/_0761_ ) );
INV_X1 \myexu/_3752_ ( .A(\myexu/_2526_ ), .ZN(\myexu/_0762_ ) );
NOR3_X1 \myexu/_3753_ ( .A1(\myexu/_0762_ ), .A2(\myexu/_2527_ ), .A3(\myexu/_2525_ ), .ZN(\myexu/_0763_ ) );
NOR2_X1 \myexu/_3754_ ( .A1(\myexu/_2118_ ), .A2(\myexu/_2524_ ), .ZN(\myexu/_0764_ ) );
AND2_X1 \myexu/_3755_ ( .A1(\myexu/_0763_ ), .A2(\myexu/_0764_ ), .ZN(\myexu/_0765_ ) );
AND2_X1 \myexu/_3756_ ( .A1(\myexu/_2527_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_0766_ ) );
NOR3_X1 \myexu/_3757_ ( .A1(fanout_net_7 ), .A2(\myexu/_2524_ ), .A3(\myexu/_2525_ ), .ZN(\myexu/_0767_ ) );
AOI21_X1 \myexu/_3758_ ( .A(\myexu/_0765_ ), .B1(\myexu/_0766_ ), .B2(\myexu/_0767_ ), .ZN(\myexu/_0768_ ) );
OR2_X1 \myexu/_3759_ ( .A1(\myexu/_0761_ ), .A2(\myexu/_0768_ ), .ZN(\myexu/_0769_ ) );
NOR2_X1 \myexu/_3760_ ( .A1(fanout_net_7 ), .A2(\myexu/_2524_ ), .ZN(\myexu/_0770_ ) );
AND2_X1 \myexu/_3761_ ( .A1(\myexu/_0763_ ), .A2(\myexu/_0770_ ), .ZN(\myexu/_0771_ ) );
INV_X1 \myexu/_3762_ ( .A(\myexu/_0771_ ), .ZN(\myexu/_0772_ ) );
BUF_X4 \myexu/_3763_ ( .A(\myexu/_0772_ ), .Z(\myexu/_0773_ ) );
XNOR2_X1 \myexu/_3764_ ( .A(\myexu/_2427_ ), .B(\myexu/_2459_ ), .ZN(\myexu/_0774_ ) );
NOR2_X1 \myexu/_3765_ ( .A1(\myexu/_0773_ ), .A2(\myexu/_0774_ ), .ZN(\myexu/_0775_ ) );
AND3_X1 \myexu/_3766_ ( .A1(\myexu/_2527_ ), .A2(\myexu/_2525_ ), .A3(\myexu/_2526_ ), .ZN(\myexu/_0776_ ) );
NOR2_X1 \myexu/_3767_ ( .A1(\myexu/_2107_ ), .A2(fanout_net_7 ), .ZN(\myexu/_0777_ ) );
AND2_X2 \myexu/_3768_ ( .A1(\myexu/_0776_ ), .A2(\myexu/_0777_ ), .ZN(\myexu/_0778_ ) );
AND2_X1 \myexu/_3769_ ( .A1(\myexu/_0776_ ), .A2(\myexu/_0770_ ), .ZN(\myexu/_0779_ ) );
BUF_X4 \myexu/_3770_ ( .A(\myexu/_0779_ ), .Z(\myexu/_0780_ ) );
XOR2_X1 \myexu/_3771_ ( .A(\myexu/_0295_ ), .B(\myexu/_2260_ ), .Z(\myexu/_0781_ ) );
AOI221_X4 \myexu/_3772_ ( .A(\myexu/_0775_ ), .B1(\myexu/_0295_ ), .B2(\myexu/_0778_ ), .C1(\myexu/_0780_ ), .C2(\myexu/_0781_ ), .ZN(\myexu/_0782_ ) );
AOI21_X1 \myexu/_3773_ ( .A(\myexu/_0640_ ), .B1(\myexu/_0769_ ), .B2(\myexu/_0782_ ), .ZN(\myexu/_0783_ ) );
AND2_X2 \myexu/_3774_ ( .A1(\myexu/_0636_ ), .A2(\myexu/_2530_ ), .ZN(\myexu/_0784_ ) );
BUF_X4 \myexu/_3775_ ( .A(\myexu/_0784_ ), .Z(\myexu/_0785_ ) );
BUF_X4 \myexu/_3776_ ( .A(\myexu/_0785_ ), .Z(\myexu/_0786_ ) );
BUF_X4 \myexu/_3777_ ( .A(\myexu/_0786_ ), .Z(\myexu/_0787_ ) );
AOI22_X1 \myexu/_3778_ ( .A1(\myexu/_0763_ ), .A2(\myexu/_0770_ ), .B1(\myexu/_0776_ ), .B2(\myexu/_2118_ ), .ZN(\myexu/_0788_ ) );
AND2_X2 \myexu/_3779_ ( .A1(\myexu/_0768_ ), .A2(\myexu/_0788_ ), .ZN(\myexu/_0789_ ) );
NOR2_X1 \myexu/_3780_ ( .A1(\myexu/_0789_ ), .A2(\myexu/_0639_ ), .ZN(\myexu/_0790_ ) );
INV_X1 \myexu/_3781_ ( .A(\myexu/_0790_ ), .ZN(\myexu/_0791_ ) );
CLKBUF_X2 \myexu/_3782_ ( .A(\myexu/_0791_ ), .Z(\myexu/_0792_ ) );
AND2_X1 \myexu/_3783_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0034_ ), .ZN(\myexu/_0793_ ) );
NOR3_X1 \myexu/_3784_ ( .A1(\myexu/_0783_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_0793_ ), .ZN(\myexu/_0794_ ) );
INV_X1 \myexu/_3785_ ( .A(\myexu/_0784_ ), .ZN(\myexu/_0795_ ) );
BUF_X4 \myexu/_3786_ ( .A(\myexu/_0795_ ), .Z(\myexu/_0796_ ) );
CLKBUF_X3 \myexu/_3787_ ( .A(\myexu/_0796_ ), .Z(\myexu/_0797_ ) );
OAI21_X1 \myexu/_3788_ ( .A(\myexu/_2156_ ), .B1(\myexu/_0797_ ), .B2(\myexu/_2260_ ), .ZN(\myexu/_0798_ ) );
OAI21_X1 \myexu/_3789_ ( .A(\myexu/_0635_ ), .B1(\myexu/_0794_ ), .B2(\myexu/_0798_ ), .ZN(\myexu/_0799_ ) );
MUX2_X1 \myexu/_3790_ ( .A(\myexu/_2394_ ), .B(\myexu/_0799_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0209_ ) );
BUF_X4 \myexu/_3791_ ( .A(\myexu/_0638_ ), .Z(\myexu/_0800_ ) );
XOR2_X2 \myexu/_3792_ ( .A(\myexu/_0306_ ), .B(\myexu/_2271_ ), .Z(\myexu/_0801_ ) );
AND2_X1 \myexu/_3793_ ( .A1(\myexu/_0295_ ), .A2(\myexu/_2260_ ), .ZN(\myexu/_0802_ ) );
XOR2_X1 \myexu/_3794_ ( .A(\myexu/_0801_ ), .B(\myexu/_0802_ ), .Z(\myexu/_0803_ ) );
INV_X1 \myexu/_3795_ ( .A(\myexu/_0803_ ), .ZN(\myexu/_0804_ ) );
INV_X1 \myexu/_3796_ ( .A(\myexu/_0779_ ), .ZN(\myexu/_0805_ ) );
INV_X1 \myexu/_3797_ ( .A(\myexu/_0778_ ), .ZN(\myexu/_0806_ ) );
OAI22_X1 \myexu/_3798_ ( .A1(\myexu/_0804_ ), .A2(\myexu/_0805_ ), .B1(\myexu/_1992_ ), .B2(\myexu/_0806_ ), .ZN(\myexu/_0807_ ) );
XNOR2_X2 \myexu/_3799_ ( .A(\myexu/_2438_ ), .B(\myexu/_2470_ ), .ZN(\myexu/_0808_ ) );
INV_X4 \myexu/_3800_ ( .A(\myexu/_0808_ ), .ZN(\myexu/_0809_ ) );
NOR2_X4 \myexu/_3801_ ( .A1(\myexu/_2103_ ), .A2(\myexu/_2427_ ), .ZN(\myexu/_0810_ ) );
OAI211_X2 \myexu/_3802_ ( .A(\myexu/_0770_ ), .B(\myexu/_0763_ ), .C1(\myexu/_0809_ ), .C2(\myexu/_0810_ ), .ZN(\myexu/_0811_ ) );
AOI21_X1 \myexu/_3803_ ( .A(\myexu/_0811_ ), .B1(\myexu/_0810_ ), .B2(\myexu/_0809_ ), .ZN(\myexu/_0812_ ) );
OAI21_X1 \myexu/_3804_ ( .A(\myexu/_0800_ ), .B1(\myexu/_0807_ ), .B2(\myexu/_0812_ ), .ZN(\myexu/_0813_ ) );
OAI21_X1 \myexu/_3805_ ( .A(\myexu/_0045_ ), .B1(\myexu/_0789_ ), .B2(\myexu/_0639_ ), .ZN(\myexu/_0814_ ) );
AOI21_X1 \myexu/_3806_ ( .A(\myexu/_0785_ ), .B1(\myexu/_0813_ ), .B2(\myexu/_0814_ ), .ZN(\myexu/_0815_ ) );
INV_X1 \myexu/_3807_ ( .A(\myexu/_2529_ ), .ZN(\myexu/_0816_ ) );
AND4_X1 \myexu/_3808_ ( .A1(\myexu/_2528_ ), .A2(\myexu/_0816_ ), .A3(\myexu/_2530_ ), .A4(\myexu/_2271_ ), .ZN(\myexu/_0817_ ) );
OR2_X1 \myexu/_3809_ ( .A1(\myexu/_0815_ ), .A2(\myexu/_0817_ ), .ZN(\myexu/_0818_ ) );
BUF_X4 \myexu/_3810_ ( .A(\myexu/_2130_ ), .Z(\myexu/_0819_ ) );
MUX2_X1 \myexu/_3811_ ( .A(\myexu/_2502_ ), .B(\myexu/_0818_ ), .S(\myexu/_0819_ ), .Z(\myexu/_0820_ ) );
MUX2_X1 \myexu/_3812_ ( .A(\myexu/_2405_ ), .B(\myexu/_0820_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0210_ ) );
NAND3_X1 \myexu/_3813_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2513_ ), .ZN(\myexu/_0821_ ) );
NAND2_X1 \myexu/_3814_ ( .A1(\myexu/_0801_ ), .A2(\myexu/_0802_ ), .ZN(\myexu/_0822_ ) );
NAND2_X1 \myexu/_3815_ ( .A1(\myexu/_0306_ ), .A2(\myexu/_2271_ ), .ZN(\myexu/_0823_ ) );
NAND2_X1 \myexu/_3816_ ( .A1(\myexu/_0822_ ), .A2(\myexu/_0823_ ), .ZN(\myexu/_0824_ ) );
XOR2_X1 \myexu/_3817_ ( .A(\myexu/_0317_ ), .B(\myexu/_2282_ ), .Z(\myexu/_0825_ ) );
XOR2_X1 \myexu/_3818_ ( .A(\myexu/_0824_ ), .B(\myexu/_0825_ ), .Z(\myexu/_0826_ ) );
BUF_X4 \myexu/_3819_ ( .A(\myexu/_0780_ ), .Z(\myexu/_0827_ ) );
BUF_X4 \myexu/_3820_ ( .A(\myexu/_0778_ ), .Z(\myexu/_0828_ ) );
AOI22_X1 \myexu/_3821_ ( .A1(\myexu/_0826_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0317_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_0829_ ) );
NAND2_X1 \myexu/_3822_ ( .A1(\myexu/_2125_ ), .A2(\myexu/_2438_ ), .ZN(\myexu/_0830_ ) );
OAI21_X4 \myexu/_3823_ ( .A(\myexu/_0830_ ), .B1(\myexu/_0809_ ), .B2(\myexu/_0810_ ), .ZN(\myexu/_0831_ ) );
XNOR2_X1 \myexu/_3824_ ( .A(\myexu/_2449_ ), .B(\myexu/_2481_ ), .ZN(\myexu/_0832_ ) );
AND2_X4 \myexu/_3825_ ( .A1(\myexu/_0831_ ), .A2(\myexu/_0832_ ), .ZN(\myexu/_0833_ ) );
BUF_X4 \myexu/_3826_ ( .A(\myexu/_0771_ ), .Z(\myexu/_0834_ ) );
OAI21_X1 \myexu/_3827_ ( .A(\myexu/_0834_ ), .B1(\myexu/_0831_ ), .B2(\myexu/_0832_ ), .ZN(\myexu/_0835_ ) );
OAI21_X1 \myexu/_3828_ ( .A(\myexu/_0829_ ), .B1(\myexu/_0833_ ), .B2(\myexu/_0835_ ), .ZN(\myexu/_0836_ ) );
NAND2_X1 \myexu/_3829_ ( .A1(\myexu/_0836_ ), .A2(\myexu/_0800_ ), .ZN(\myexu/_0837_ ) );
OAI21_X1 \myexu/_3830_ ( .A(\myexu/_0056_ ), .B1(\myexu/_0789_ ), .B2(\myexu/_0639_ ), .ZN(\myexu/_0838_ ) );
AND3_X1 \myexu/_3831_ ( .A1(\myexu/_0837_ ), .A2(\myexu/_0796_ ), .A3(\myexu/_0838_ ), .ZN(\myexu/_0839_ ) );
INV_X1 \myexu/_3832_ ( .A(\myexu/_2282_ ), .ZN(\myexu/_0840_ ) );
OAI21_X1 \myexu/_3833_ ( .A(\myexu/_2156_ ), .B1(\myexu/_0797_ ), .B2(\myexu/_0840_ ), .ZN(\myexu/_0841_ ) );
OAI21_X1 \myexu/_3834_ ( .A(\myexu/_0821_ ), .B1(\myexu/_0839_ ), .B2(\myexu/_0841_ ), .ZN(\myexu/_0842_ ) );
MUX2_X1 \myexu/_3835_ ( .A(\myexu/_2416_ ), .B(\myexu/_0842_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0211_ ) );
OAI21_X1 \myexu/_3836_ ( .A(\myexu/_2419_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_0843_ ) );
NAND2_X2 \myexu/_3837_ ( .A1(\myexu/_1975_ ), .A2(\myexu/_2049_ ), .ZN(\myexu/_0844_ ) );
BUF_X4 \myexu/_3838_ ( .A(\myexu/_0639_ ), .Z(\myexu/_0845_ ) );
NAND2_X1 \myexu/_3839_ ( .A1(\myexu/_0824_ ), .A2(\myexu/_0825_ ), .ZN(\myexu/_0846_ ) );
AND2_X1 \myexu/_3840_ ( .A1(\myexu/_0317_ ), .A2(\myexu/_2282_ ), .ZN(\myexu/_0847_ ) );
INV_X1 \myexu/_3841_ ( .A(\myexu/_0847_ ), .ZN(\myexu/_0848_ ) );
NAND2_X1 \myexu/_3842_ ( .A1(\myexu/_0846_ ), .A2(\myexu/_0848_ ), .ZN(\myexu/_0849_ ) );
XOR2_X1 \myexu/_3843_ ( .A(\myexu/_0320_ ), .B(\myexu/_2285_ ), .Z(\myexu/_0850_ ) );
XNOR2_X1 \myexu/_3844_ ( .A(\myexu/_0849_ ), .B(\myexu/_0850_ ), .ZN(\myexu/_0851_ ) );
INV_X1 \myexu/_3845_ ( .A(\myexu/_0851_ ), .ZN(\myexu/_0852_ ) );
BUF_X4 \myexu/_3846_ ( .A(\myexu/_0780_ ), .Z(\myexu/_0853_ ) );
BUF_X4 \myexu/_3847_ ( .A(\myexu/_0778_ ), .Z(\myexu/_0854_ ) );
AOI22_X1 \myexu/_3848_ ( .A1(\myexu/_0852_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0320_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_0855_ ) );
NOR2_X1 \myexu/_3849_ ( .A1(\myexu/_2137_ ), .A2(\myexu/_2481_ ), .ZN(\myexu/_0856_ ) );
XNOR2_X1 \myexu/_3850_ ( .A(\myexu/_2452_ ), .B(\myexu/_2484_ ), .ZN(\myexu/_0857_ ) );
OR3_X1 \myexu/_3851_ ( .A1(\myexu/_0833_ ), .A2(\myexu/_0856_ ), .A3(\myexu/_0857_ ), .ZN(\myexu/_0858_ ) );
OAI21_X4 \myexu/_3852_ ( .A(\myexu/_0857_ ), .B1(\myexu/_0833_ ), .B2(\myexu/_0856_ ), .ZN(\myexu/_0859_ ) );
NAND3_X1 \myexu/_3853_ ( .A1(\myexu/_0858_ ), .A2(\myexu/_0834_ ), .A3(\myexu/_0859_ ), .ZN(\myexu/_0860_ ) );
AOI21_X1 \myexu/_3854_ ( .A(\myexu/_0845_ ), .B1(\myexu/_0855_ ), .B2(\myexu/_0860_ ), .ZN(\myexu/_0861_ ) );
BUF_X4 \myexu/_3855_ ( .A(\myexu/_0787_ ), .Z(\myexu/_0862_ ) );
AND2_X1 \myexu/_3856_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0059_ ), .ZN(\myexu/_0863_ ) );
NOR3_X1 \myexu/_3857_ ( .A1(\myexu/_0861_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_0863_ ), .ZN(\myexu/_0864_ ) );
BUF_X4 \myexu/_3858_ ( .A(\myexu/_0796_ ), .Z(\myexu/_0865_ ) );
BUF_X4 \myexu/_3859_ ( .A(\myexu/_0865_ ), .Z(\myexu/_0866_ ) );
XOR2_X1 \myexu/_3860_ ( .A(\myexu/_2282_ ), .B(\myexu/_2285_ ), .Z(\myexu/_0867_ ) );
OAI211_X2 \myexu/_3861_ ( .A(\myexu/_1976_ ), .B(\myexu/_2140_ ), .C1(\myexu/_0866_ ), .C2(\myexu/_0867_ ), .ZN(\myexu/_0868_ ) );
OAI221_X1 \myexu/_3862_ ( .A(\myexu/_0843_ ), .B1(\myexu/_2146_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_0864_ ), .C2(\myexu/_0868_ ), .ZN(\myexu/_0212_ ) );
NAND3_X1 \myexu/_3863_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2517_ ), .ZN(\myexu/_0869_ ) );
AOI22_X1 \myexu/_3864_ ( .A1(\myexu/_0846_ ), .A2(\myexu/_0848_ ), .B1(\myexu/_1931_ ), .B2(\myexu/_2150_ ), .ZN(\myexu/_0870_ ) );
AND2_X1 \myexu/_3865_ ( .A1(\myexu/_0320_ ), .A2(\myexu/_2285_ ), .ZN(\myexu/_0871_ ) );
OR2_X1 \myexu/_3866_ ( .A1(\myexu/_0870_ ), .A2(\myexu/_0871_ ), .ZN(\myexu/_0872_ ) );
XOR2_X1 \myexu/_3867_ ( .A(\myexu/_0321_ ), .B(\myexu/_2286_ ), .Z(\myexu/_0873_ ) );
INV_X1 \myexu/_3868_ ( .A(\myexu/_0873_ ), .ZN(\myexu/_0874_ ) );
XNOR2_X1 \myexu/_3869_ ( .A(\myexu/_0872_ ), .B(\myexu/_0874_ ), .ZN(\myexu/_0875_ ) );
AOI22_X1 \myexu/_3870_ ( .A1(\myexu/_0875_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0321_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_0876_ ) );
NOR2_X1 \myexu/_3871_ ( .A1(\myexu/_0668_ ), .A2(\myexu/_2484_ ), .ZN(\myexu/_0877_ ) );
INV_X1 \myexu/_3872_ ( .A(\myexu/_0877_ ), .ZN(\myexu/_0878_ ) );
AND2_X4 \myexu/_3873_ ( .A1(\myexu/_0859_ ), .A2(\myexu/_0878_ ), .ZN(\myexu/_0879_ ) );
XNOR2_X1 \myexu/_3874_ ( .A(\myexu/_2453_ ), .B(\myexu/_2485_ ), .ZN(\myexu/_0880_ ) );
INV_X1 \myexu/_3875_ ( .A(\myexu/_0880_ ), .ZN(\myexu/_0881_ ) );
AOI21_X1 \myexu/_3876_ ( .A(\myexu/_0773_ ), .B1(\myexu/_0879_ ), .B2(\myexu/_0881_ ), .ZN(\myexu/_0882_ ) );
OAI21_X1 \myexu/_3877_ ( .A(\myexu/_0882_ ), .B1(\myexu/_0879_ ), .B2(\myexu/_0881_ ), .ZN(\myexu/_0883_ ) );
AOI21_X1 \myexu/_3878_ ( .A(\myexu/_0640_ ), .B1(\myexu/_0876_ ), .B2(\myexu/_0883_ ), .ZN(\myexu/_0884_ ) );
CLKBUF_X2 \myexu/_3879_ ( .A(\myexu/_0791_ ), .Z(\myexu/_0885_ ) );
AND2_X1 \myexu/_3880_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0060_ ), .ZN(\myexu/_0886_ ) );
NOR3_X1 \myexu/_3881_ ( .A1(\myexu/_0884_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_0886_ ), .ZN(\myexu/_0887_ ) );
AND2_X4 \myexu/_3882_ ( .A1(\myexu/_2282_ ), .A2(\myexu/_2285_ ), .ZN(\myexu/_0888_ ) );
INV_X1 \myexu/_3883_ ( .A(\myexu/_2286_ ), .ZN(\myexu/_0889_ ) );
XNOR2_X1 \myexu/_3884_ ( .A(\myexu/_0888_ ), .B(\myexu/_0889_ ), .ZN(\myexu/_0890_ ) );
OAI21_X1 \myexu/_3885_ ( .A(\myexu/_2156_ ), .B1(\myexu/_0865_ ), .B2(\myexu/_0890_ ), .ZN(\myexu/_0891_ ) );
OAI21_X1 \myexu/_3886_ ( .A(\myexu/_0869_ ), .B1(\myexu/_0887_ ), .B2(\myexu/_0891_ ), .ZN(\myexu/_0892_ ) );
MUX2_X1 \myexu/_3887_ ( .A(\myexu/_2420_ ), .B(\myexu/_0892_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0213_ ) );
XNOR2_X1 \myexu/_3888_ ( .A(\myexu/_2454_ ), .B(\myexu/_2486_ ), .ZN(\myexu/_0893_ ) );
NOR2_X4 \myexu/_3889_ ( .A1(\myexu/_0879_ ), .A2(\myexu/_0881_ ), .ZN(\myexu/_0894_ ) );
NOR2_X1 \myexu/_3890_ ( .A1(\myexu/_0682_ ), .A2(\myexu/_2485_ ), .ZN(\myexu/_0895_ ) );
OAI21_X2 \myexu/_3891_ ( .A(\myexu/_0893_ ), .B1(\myexu/_0894_ ), .B2(\myexu/_0895_ ), .ZN(\myexu/_0896_ ) );
INV_X2 \myexu/_3892_ ( .A(\myexu/_0896_ ), .ZN(\myexu/_0897_ ) );
NOR3_X1 \myexu/_3893_ ( .A1(\myexu/_0894_ ), .A2(\myexu/_0895_ ), .A3(\myexu/_0893_ ), .ZN(\myexu/_0898_ ) );
NOR3_X1 \myexu/_3894_ ( .A1(\myexu/_0897_ ), .A2(\myexu/_0898_ ), .A3(\myexu/_0773_ ), .ZN(\myexu/_0899_ ) );
OAI21_X1 \myexu/_3895_ ( .A(\myexu/_0873_ ), .B1(\myexu/_0870_ ), .B2(\myexu/_0871_ ), .ZN(\myexu/_0900_ ) );
NAND2_X1 \myexu/_3896_ ( .A1(\myexu/_0321_ ), .A2(\myexu/_2286_ ), .ZN(\myexu/_0901_ ) );
NAND2_X1 \myexu/_3897_ ( .A1(\myexu/_0900_ ), .A2(\myexu/_0901_ ), .ZN(\myexu/_0902_ ) );
XOR2_X1 \myexu/_3898_ ( .A(\myexu/_0322_ ), .B(\myexu/_2287_ ), .Z(\myexu/_0903_ ) );
XNOR2_X1 \myexu/_3899_ ( .A(\myexu/_0902_ ), .B(\myexu/_0903_ ), .ZN(\myexu/_0904_ ) );
OAI22_X1 \myexu/_3900_ ( .A1(\myexu/_0904_ ), .A2(\myexu/_0805_ ), .B1(\myexu/_2164_ ), .B2(\myexu/_0806_ ), .ZN(\myexu/_0905_ ) );
OAI21_X1 \myexu/_3901_ ( .A(\myexu/_0800_ ), .B1(\myexu/_0899_ ), .B2(\myexu/_0905_ ), .ZN(\myexu/_0906_ ) );
AOI21_X1 \myexu/_3902_ ( .A(\myexu/_0785_ ), .B1(\myexu/_0791_ ), .B2(\myexu/_0061_ ), .ZN(\myexu/_0907_ ) );
AND2_X4 \myexu/_3903_ ( .A1(\myexu/_0888_ ), .A2(\myexu/_2286_ ), .ZN(\myexu/_0908_ ) );
XNOR2_X1 \myexu/_3904_ ( .A(\myexu/_0908_ ), .B(\myexu/_2287_ ), .ZN(\myexu/_0909_ ) );
AOI22_X1 \myexu/_3905_ ( .A1(\myexu/_0906_ ), .A2(\myexu/_0907_ ), .B1(\myexu/_0786_ ), .B2(\myexu/_0909_ ), .ZN(\myexu/_0910_ ) );
MUX2_X1 \myexu/_3906_ ( .A(\myexu/_2518_ ), .B(\myexu/_0910_ ), .S(\myexu/_2131_ ), .Z(\myexu/_0911_ ) );
MUX2_X1 \myexu/_3907_ ( .A(\myexu/_2421_ ), .B(\myexu/_0911_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0214_ ) );
OAI21_X1 \myexu/_3908_ ( .A(\myexu/_2422_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_0912_ ) );
BUF_X4 \myexu/_3909_ ( .A(\myexu/_0773_ ), .Z(\myexu/_0913_ ) );
INV_X1 \myexu/_3910_ ( .A(\myexu/_2486_ ), .ZN(\myexu/_0914_ ) );
AOI21_X4 \myexu/_3911_ ( .A(\myexu/_0897_ ), .B1(\myexu/_2454_ ), .B2(\myexu/_0914_ ), .ZN(\myexu/_0915_ ) );
XNOR2_X1 \myexu/_3912_ ( .A(\myexu/_2455_ ), .B(\myexu/_2487_ ), .ZN(\myexu/_0916_ ) );
INV_X1 \myexu/_3913_ ( .A(\myexu/_0916_ ), .ZN(\myexu/_0917_ ) );
AOI21_X1 \myexu/_3914_ ( .A(\myexu/_0913_ ), .B1(\myexu/_0915_ ), .B2(\myexu/_0917_ ), .ZN(\myexu/_0918_ ) );
OAI21_X1 \myexu/_3915_ ( .A(\myexu/_0918_ ), .B1(\myexu/_0915_ ), .B2(\myexu/_0917_ ), .ZN(\myexu/_0919_ ) );
AND3_X1 \myexu/_3916_ ( .A1(\myexu/_0903_ ), .A2(\myexu/_0321_ ), .A3(\myexu/_2286_ ), .ZN(\myexu/_0920_ ) );
AND2_X1 \myexu/_3917_ ( .A1(\myexu/_0322_ ), .A2(\myexu/_2287_ ), .ZN(\myexu/_0921_ ) );
OR2_X1 \myexu/_3918_ ( .A1(\myexu/_0920_ ), .A2(\myexu/_0921_ ), .ZN(\myexu/_0922_ ) );
AND2_X1 \myexu/_3919_ ( .A1(\myexu/_0873_ ), .A2(\myexu/_0903_ ), .ZN(\myexu/_0923_ ) );
AOI21_X1 \myexu/_3920_ ( .A(\myexu/_0922_ ), .B1(\myexu/_0872_ ), .B2(\myexu/_0923_ ), .ZN(\myexu/_0924_ ) );
XOR2_X1 \myexu/_3921_ ( .A(\myexu/_0323_ ), .B(\myexu/_2288_ ), .Z(\myexu/_0925_ ) );
XNOR2_X1 \myexu/_3922_ ( .A(\myexu/_0924_ ), .B(\myexu/_0925_ ), .ZN(\myexu/_0926_ ) );
AOI22_X1 \myexu/_3923_ ( .A1(\myexu/_0926_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0323_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_0927_ ) );
AOI21_X1 \myexu/_3924_ ( .A(\myexu/_0845_ ), .B1(\myexu/_0919_ ), .B2(\myexu/_0927_ ), .ZN(\myexu/_0928_ ) );
AND2_X1 \myexu/_3925_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0062_ ), .ZN(\myexu/_0929_ ) );
NOR3_X1 \myexu/_3926_ ( .A1(\myexu/_0928_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_0929_ ), .ZN(\myexu/_0930_ ) );
AND2_X2 \myexu/_3927_ ( .A1(\myexu/_0819_ ), .A2(\myexu/_1974_ ), .ZN(\myexu/_0931_ ) );
AND2_X1 \myexu/_3928_ ( .A1(\myexu/_0908_ ), .A2(\myexu/_2287_ ), .ZN(\myexu/_0932_ ) );
XNOR2_X1 \myexu/_3929_ ( .A(\myexu/_0932_ ), .B(\myexu/_2177_ ), .ZN(\myexu/_0933_ ) );
OAI21_X1 \myexu/_3930_ ( .A(\myexu/_0931_ ), .B1(\myexu/_0933_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_0934_ ) );
OAI221_X1 \myexu/_3931_ ( .A(\myexu/_0912_ ), .B1(\myexu/_2172_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_0930_ ), .C2(\myexu/_0934_ ), .ZN(\myexu/_0215_ ) );
NAND3_X1 \myexu/_3932_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2520_ ), .ZN(\myexu/_0935_ ) );
NOR2_X1 \myexu/_3933_ ( .A1(\myexu/_0323_ ), .A2(\myexu/_2288_ ), .ZN(\myexu/_0936_ ) );
AND2_X1 \myexu/_3934_ ( .A1(\myexu/_0323_ ), .A2(\myexu/_2288_ ), .ZN(\myexu/_0937_ ) );
NOR3_X1 \myexu/_3935_ ( .A1(\myexu/_0924_ ), .A2(\myexu/_0936_ ), .A3(\myexu/_0937_ ), .ZN(\myexu/_0938_ ) );
NOR2_X1 \myexu/_3936_ ( .A1(\myexu/_0938_ ), .A2(\myexu/_0937_ ), .ZN(\myexu/_0939_ ) );
XOR2_X1 \myexu/_3937_ ( .A(\myexu/_0324_ ), .B(\myexu/_2289_ ), .Z(\myexu/_0940_ ) );
XNOR2_X1 \myexu/_3938_ ( .A(\myexu/_0939_ ), .B(\myexu/_0940_ ), .ZN(\myexu/_0941_ ) );
AOI22_X1 \myexu/_3939_ ( .A1(\myexu/_0941_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0324_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_0942_ ) );
NOR2_X4 \myexu/_3940_ ( .A1(\myexu/_0915_ ), .A2(\myexu/_0917_ ), .ZN(\myexu/_0943_ ) );
AOI21_X4 \myexu/_3941_ ( .A(\myexu/_0943_ ), .B1(\myexu/_2455_ ), .B2(\myexu/_2176_ ), .ZN(\myexu/_0944_ ) );
XNOR2_X1 \myexu/_3942_ ( .A(\myexu/_2456_ ), .B(\myexu/_2488_ ), .ZN(\myexu/_0945_ ) );
XOR2_X1 \myexu/_3943_ ( .A(\myexu/_0944_ ), .B(\myexu/_0945_ ), .Z(\myexu/_0946_ ) );
OAI21_X1 \myexu/_3944_ ( .A(\myexu/_0942_ ), .B1(\myexu/_0946_ ), .B2(\myexu/_0913_ ), .ZN(\myexu/_0947_ ) );
NAND2_X1 \myexu/_3945_ ( .A1(\myexu/_0947_ ), .A2(\myexu/_0800_ ), .ZN(\myexu/_0948_ ) );
OAI21_X1 \myexu/_3946_ ( .A(\myexu/_0063_ ), .B1(\myexu/_0789_ ), .B2(\myexu/_0639_ ), .ZN(\myexu/_0949_ ) );
AND3_X1 \myexu/_3947_ ( .A1(\myexu/_0948_ ), .A2(\myexu/_0796_ ), .A3(\myexu/_0949_ ), .ZN(\myexu/_0950_ ) );
AND2_X1 \myexu/_3948_ ( .A1(\myexu/_0932_ ), .A2(\myexu/_2288_ ), .ZN(\myexu/_0951_ ) );
INV_X1 \myexu/_3949_ ( .A(\myexu/_2289_ ), .ZN(\myexu/_0952_ ) );
XNOR2_X1 \myexu/_3950_ ( .A(\myexu/_0951_ ), .B(\myexu/_0952_ ), .ZN(\myexu/_0953_ ) );
OAI21_X1 \myexu/_3951_ ( .A(\myexu/_2156_ ), .B1(\myexu/_0953_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_0954_ ) );
OAI21_X1 \myexu/_3952_ ( .A(\myexu/_0935_ ), .B1(\myexu/_0950_ ), .B2(\myexu/_0954_ ), .ZN(\myexu/_0955_ ) );
MUX2_X1 \myexu/_3953_ ( .A(\myexu/_2423_ ), .B(\myexu/_0955_ ), .S(\myexu/_0616_ ), .Z(\myexu/_0216_ ) );
NAND3_X1 \myexu/_3954_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2521_ ), .ZN(\myexu/_0956_ ) );
AOI21_X4 \myexu/_3955_ ( .A(\myexu/_0944_ ), .B1(\myexu/_2181_ ), .B2(\myexu/_2488_ ), .ZN(\myexu/_0957_ ) );
NOR2_X1 \myexu/_3956_ ( .A1(\myexu/_2181_ ), .A2(\myexu/_2488_ ), .ZN(\myexu/_0958_ ) );
NOR2_X4 \myexu/_3957_ ( .A1(\myexu/_0957_ ), .A2(\myexu/_0958_ ), .ZN(\myexu/_0959_ ) );
INV_X4 \myexu/_3958_ ( .A(\myexu/_0959_ ), .ZN(\myexu/_0960_ ) );
XNOR2_X1 \myexu/_3959_ ( .A(\myexu/_2457_ ), .B(\myexu/_2489_ ), .ZN(\myexu/_0961_ ) );
AND2_X1 \myexu/_3960_ ( .A1(\myexu/_0960_ ), .A2(\myexu/_0961_ ), .ZN(\myexu/_0962_ ) );
NOR3_X1 \myexu/_3961_ ( .A1(\myexu/_0957_ ), .A2(\myexu/_0958_ ), .A3(\myexu/_0961_ ), .ZN(\myexu/_0963_ ) );
OR3_X1 \myexu/_3962_ ( .A1(\myexu/_0962_ ), .A2(\myexu/_0773_ ), .A3(\myexu/_0963_ ), .ZN(\myexu/_0964_ ) );
AND2_X1 \myexu/_3963_ ( .A1(\myexu/_0925_ ), .A2(\myexu/_0940_ ), .ZN(\myexu/_0965_ ) );
OAI211_X2 \myexu/_3964_ ( .A(\myexu/_0923_ ), .B(\myexu/_0965_ ), .C1(\myexu/_0870_ ), .C2(\myexu/_0871_ ), .ZN(\myexu/_0966_ ) );
AND2_X1 \myexu/_3965_ ( .A1(\myexu/_0940_ ), .A2(\myexu/_0937_ ), .ZN(\myexu/_0967_ ) );
AOI221_X4 \myexu/_3966_ ( .A(\myexu/_0967_ ), .B1(\myexu/_0324_ ), .B2(\myexu/_2289_ ), .C1(\myexu/_0922_ ), .C2(\myexu/_0965_ ), .ZN(\myexu/_0968_ ) );
NAND2_X4 \myexu/_3967_ ( .A1(\myexu/_0966_ ), .A2(\myexu/_0968_ ), .ZN(\myexu/_0969_ ) );
XOR2_X1 \myexu/_3968_ ( .A(\myexu/_0325_ ), .B(\myexu/_2290_ ), .Z(\myexu/_0970_ ) );
XOR2_X1 \myexu/_3969_ ( .A(\myexu/_0969_ ), .B(\myexu/_0970_ ), .Z(\myexu/_0971_ ) );
AOI22_X1 \myexu/_3970_ ( .A1(\myexu/_0971_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0325_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_0972_ ) );
AOI21_X1 \myexu/_3971_ ( .A(\myexu/_0640_ ), .B1(\myexu/_0964_ ), .B2(\myexu/_0972_ ), .ZN(\myexu/_0973_ ) );
AND2_X1 \myexu/_3972_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0064_ ), .ZN(\myexu/_0974_ ) );
NOR3_X1 \myexu/_3973_ ( .A1(\myexu/_0973_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_0974_ ), .ZN(\myexu/_0975_ ) );
AND2_X2 \myexu/_3974_ ( .A1(\myexu/_0951_ ), .A2(\myexu/_2289_ ), .ZN(\myexu/_0976_ ) );
INV_X1 \myexu/_3975_ ( .A(\myexu/_2290_ ), .ZN(\myexu/_0977_ ) );
XNOR2_X1 \myexu/_3976_ ( .A(\myexu/_0976_ ), .B(\myexu/_0977_ ), .ZN(\myexu/_0978_ ) );
OAI21_X1 \myexu/_3977_ ( .A(\myexu/_0819_ ), .B1(\myexu/_0978_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_0979_ ) );
OAI21_X1 \myexu/_3978_ ( .A(\myexu/_0956_ ), .B1(\myexu/_0975_ ), .B2(\myexu/_0979_ ), .ZN(\myexu/_0980_ ) );
BUF_X4 \myexu/_3979_ ( .A(\myexu/_1974_ ), .Z(\myexu/_0981_ ) );
MUX2_X1 \myexu/_3980_ ( .A(\myexu/_2424_ ), .B(\myexu/_0980_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0217_ ) );
OAI21_X1 \myexu/_3981_ ( .A(\myexu/_2425_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_0982_ ) );
NOR2_X1 \myexu/_3982_ ( .A1(\myexu/_0697_ ), .A2(\myexu/_2489_ ), .ZN(\myexu/_0983_ ) );
XNOR2_X1 \myexu/_3983_ ( .A(\myexu/_2458_ ), .B(\myexu/_2490_ ), .ZN(\myexu/_0984_ ) );
NOR3_X1 \myexu/_3984_ ( .A1(\myexu/_0962_ ), .A2(\myexu/_0983_ ), .A3(\myexu/_0984_ ), .ZN(\myexu/_0985_ ) );
AND2_X1 \myexu/_3985_ ( .A1(\myexu/_0984_ ), .A2(\myexu/_0983_ ), .ZN(\myexu/_0986_ ) );
NOR2_X1 \myexu/_3986_ ( .A1(\myexu/_0913_ ), .A2(\myexu/_0986_ ), .ZN(\myexu/_0987_ ) );
NAND2_X1 \myexu/_3987_ ( .A1(\myexu/_0961_ ), .A2(\myexu/_0984_ ), .ZN(\myexu/_0988_ ) );
OAI21_X1 \myexu/_3988_ ( .A(\myexu/_0987_ ), .B1(\myexu/_0959_ ), .B2(\myexu/_0988_ ), .ZN(\myexu/_0989_ ) );
NOR2_X1 \myexu/_3989_ ( .A1(\myexu/_0985_ ), .A2(\myexu/_0989_ ), .ZN(\myexu/_0990_ ) );
NAND3_X1 \myexu/_3990_ ( .A1(\myexu/_0776_ ), .A2(\myexu/_0777_ ), .A3(\myexu/_0326_ ), .ZN(\myexu/_0991_ ) );
NAND2_X1 \myexu/_3991_ ( .A1(\myexu/_0969_ ), .A2(\myexu/_0970_ ), .ZN(\myexu/_0992_ ) );
NAND2_X1 \myexu/_3992_ ( .A1(\myexu/_0325_ ), .A2(\myexu/_2290_ ), .ZN(\myexu/_0993_ ) );
NAND2_X1 \myexu/_3993_ ( .A1(\myexu/_0992_ ), .A2(\myexu/_0993_ ), .ZN(\myexu/_0994_ ) );
AND2_X1 \myexu/_3994_ ( .A1(\myexu/_0326_ ), .A2(\myexu/_2291_ ), .ZN(\myexu/_0995_ ) );
NOR2_X1 \myexu/_3995_ ( .A1(\myexu/_0326_ ), .A2(\myexu/_2291_ ), .ZN(\myexu/_0996_ ) );
NOR2_X1 \myexu/_3996_ ( .A1(\myexu/_0995_ ), .A2(\myexu/_0996_ ), .ZN(\myexu/_0997_ ) );
XNOR2_X1 \myexu/_3997_ ( .A(\myexu/_0994_ ), .B(\myexu/_0997_ ), .ZN(\myexu/_0998_ ) );
OAI21_X1 \myexu/_3998_ ( .A(\myexu/_0991_ ), .B1(\myexu/_0998_ ), .B2(\myexu/_0805_ ), .ZN(\myexu/_0999_ ) );
OAI21_X1 \myexu/_3999_ ( .A(\myexu/_0800_ ), .B1(\myexu/_0990_ ), .B2(\myexu/_0999_ ), .ZN(\myexu/_1000_ ) );
OAI21_X1 \myexu/_4000_ ( .A(\myexu/_0065_ ), .B1(\myexu/_0789_ ), .B2(\myexu/_0845_ ), .ZN(\myexu/_1001_ ) );
AND3_X1 \myexu/_4001_ ( .A1(\myexu/_1000_ ), .A2(\myexu/_0866_ ), .A3(\myexu/_1001_ ), .ZN(\myexu/_1002_ ) );
AND2_X2 \myexu/_4002_ ( .A1(\myexu/_0976_ ), .A2(\myexu/_2290_ ), .ZN(\myexu/_1003_ ) );
XNOR2_X1 \myexu/_4003_ ( .A(\myexu/_1003_ ), .B(\myexu/_2291_ ), .ZN(\myexu/_1004_ ) );
NAND2_X1 \myexu/_4004_ ( .A1(\myexu/_1004_ ), .A2(\myexu/_0862_ ), .ZN(\myexu/_1005_ ) );
NAND2_X1 \myexu/_4005_ ( .A1(\myexu/_1005_ ), .A2(\myexu/_0931_ ), .ZN(\myexu/_1006_ ) );
OAI221_X1 \myexu/_4006_ ( .A(\myexu/_0982_ ), .B1(\myexu/_2198_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1002_ ), .C2(\myexu/_1006_ ), .ZN(\myexu/_0218_ ) );
OAI21_X1 \myexu/_4007_ ( .A(\myexu/_2395_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1007_ ) );
AOI21_X1 \myexu/_4008_ ( .A(\myexu/_0986_ ), .B1(\myexu/_2458_ ), .B2(\myexu/_2202_ ), .ZN(\myexu/_1008_ ) );
OAI21_X1 \myexu/_4009_ ( .A(\myexu/_1008_ ), .B1(\myexu/_0959_ ), .B2(\myexu/_0988_ ), .ZN(\myexu/_1009_ ) );
XNOR2_X1 \myexu/_4010_ ( .A(\myexu/_2428_ ), .B(\myexu/_2460_ ), .ZN(\myexu/_1010_ ) );
AND2_X1 \myexu/_4011_ ( .A1(\myexu/_1009_ ), .A2(\myexu/_1010_ ), .ZN(\myexu/_1011_ ) );
OAI21_X1 \myexu/_4012_ ( .A(\myexu/_0834_ ), .B1(\myexu/_1009_ ), .B2(\myexu/_1010_ ), .ZN(\myexu/_1012_ ) );
OR2_X1 \myexu/_4013_ ( .A1(\myexu/_1011_ ), .A2(\myexu/_1012_ ), .ZN(\myexu/_1013_ ) );
NOR3_X1 \myexu/_4014_ ( .A1(\myexu/_0995_ ), .A2(\myexu/_0996_ ), .A3(\myexu/_0993_ ), .ZN(\myexu/_1014_ ) );
OR2_X1 \myexu/_4015_ ( .A1(\myexu/_1014_ ), .A2(\myexu/_0995_ ), .ZN(\myexu/_1015_ ) );
AND2_X1 \myexu/_4016_ ( .A1(\myexu/_0970_ ), .A2(\myexu/_0997_ ), .ZN(\myexu/_1016_ ) );
AOI21_X1 \myexu/_4017_ ( .A(\myexu/_1015_ ), .B1(\myexu/_0969_ ), .B2(\myexu/_1016_ ), .ZN(\myexu/_1017_ ) );
XNOR2_X1 \myexu/_4018_ ( .A(\myexu/_0296_ ), .B(\myexu/_2261_ ), .ZN(\myexu/_1018_ ) );
XOR2_X1 \myexu/_4019_ ( .A(\myexu/_1017_ ), .B(\myexu/_1018_ ), .Z(\myexu/_1019_ ) );
AOI22_X1 \myexu/_4020_ ( .A1(\myexu/_1019_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0296_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1020_ ) );
AOI21_X1 \myexu/_4021_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1013_ ), .B2(\myexu/_1020_ ), .ZN(\myexu/_1021_ ) );
AND2_X1 \myexu/_4022_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0035_ ), .ZN(\myexu/_1022_ ) );
NOR3_X1 \myexu/_4023_ ( .A1(\myexu/_1021_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1022_ ), .ZN(\myexu/_1023_ ) );
AND2_X4 \myexu/_4024_ ( .A1(\myexu/_1003_ ), .A2(\myexu/_2291_ ), .ZN(\myexu/_1024_ ) );
INV_X1 \myexu/_4025_ ( .A(\myexu/_2261_ ), .ZN(\myexu/_1025_ ) );
XNOR2_X1 \myexu/_4026_ ( .A(\myexu/_1024_ ), .B(\myexu/_1025_ ), .ZN(\myexu/_1026_ ) );
OAI21_X1 \myexu/_4027_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1026_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1027_ ) );
OAI221_X1 \myexu/_4028_ ( .A(\myexu/_1007_ ), .B1(\myexu/_2211_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1023_ ), .C2(\myexu/_1027_ ), .ZN(\myexu/_0219_ ) );
INV_X1 \myexu/_4029_ ( .A(\myexu/_2216_ ), .ZN(\myexu/_1028_ ) );
NOR2_X1 \myexu/_4030_ ( .A1(\myexu/_2210_ ), .A2(\myexu/_2460_ ), .ZN(\myexu/_1029_ ) );
XNOR2_X1 \myexu/_4031_ ( .A(\myexu/_2429_ ), .B(\myexu/_2461_ ), .ZN(\myexu/_1030_ ) );
OR3_X1 \myexu/_4032_ ( .A1(\myexu/_1011_ ), .A2(\myexu/_1029_ ), .A3(\myexu/_1030_ ), .ZN(\myexu/_1031_ ) );
OAI21_X1 \myexu/_4033_ ( .A(\myexu/_1030_ ), .B1(\myexu/_1011_ ), .B2(\myexu/_1029_ ), .ZN(\myexu/_1032_ ) );
NAND3_X1 \myexu/_4034_ ( .A1(\myexu/_1031_ ), .A2(\myexu/_0834_ ), .A3(\myexu/_1032_ ), .ZN(\myexu/_1033_ ) );
NOR2_X1 \myexu/_4035_ ( .A1(\myexu/_1017_ ), .A2(\myexu/_1018_ ), .ZN(\myexu/_1034_ ) );
AND2_X1 \myexu/_4036_ ( .A1(\myexu/_0296_ ), .A2(\myexu/_2261_ ), .ZN(\myexu/_1035_ ) );
NOR2_X1 \myexu/_4037_ ( .A1(\myexu/_1034_ ), .A2(\myexu/_1035_ ), .ZN(\myexu/_1036_ ) );
XOR2_X1 \myexu/_4038_ ( .A(\myexu/_0297_ ), .B(\myexu/_2262_ ), .Z(\myexu/_1037_ ) );
XNOR2_X1 \myexu/_4039_ ( .A(\myexu/_1036_ ), .B(\myexu/_1037_ ), .ZN(\myexu/_1038_ ) );
AOI22_X1 \myexu/_4040_ ( .A1(\myexu/_1038_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0297_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1039_ ) );
AOI21_X1 \myexu/_4041_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1033_ ), .B2(\myexu/_1039_ ), .ZN(\myexu/_1040_ ) );
AND2_X1 \myexu/_4042_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0036_ ), .ZN(\myexu/_1041_ ) );
NOR3_X1 \myexu/_4043_ ( .A1(\myexu/_1040_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_1041_ ), .ZN(\myexu/_1042_ ) );
AND2_X1 \myexu/_4044_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_2261_ ), .ZN(\myexu/_1043_ ) );
XOR2_X1 \myexu/_4045_ ( .A(\myexu/_1043_ ), .B(\myexu/_2262_ ), .Z(\myexu/_1044_ ) );
OAI21_X1 \myexu/_4046_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1044_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_1045_ ) );
OAI21_X1 \myexu/_4047_ ( .A(\myexu/_1028_ ), .B1(\myexu/_1042_ ), .B2(\myexu/_1045_ ), .ZN(\myexu/_1046_ ) );
MUX2_X1 \myexu/_4048_ ( .A(\myexu/_2396_ ), .B(\myexu/_1046_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0220_ ) );
OAI21_X1 \myexu/_4049_ ( .A(\myexu/_2397_ ), .B1(\myexu/_1983_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1047_ ) );
NAND2_X1 \myexu/_4050_ ( .A1(\myexu/_1010_ ), .A2(\myexu/_1030_ ), .ZN(\myexu/_1048_ ) );
NOR2_X1 \myexu/_4051_ ( .A1(\myexu/_1008_ ), .A2(\myexu/_1048_ ), .ZN(\myexu/_1049_ ) );
NOR2_X1 \myexu/_4052_ ( .A1(\myexu/_0700_ ), .A2(\myexu/_2461_ ), .ZN(\myexu/_1050_ ) );
AND2_X1 \myexu/_4053_ ( .A1(\myexu/_1030_ ), .A2(\myexu/_1029_ ), .ZN(\myexu/_1051_ ) );
OR3_X1 \myexu/_4054_ ( .A1(\myexu/_1049_ ), .A2(\myexu/_1050_ ), .A3(\myexu/_1051_ ), .ZN(\myexu/_1052_ ) );
NOR2_X1 \myexu/_4055_ ( .A1(\myexu/_0988_ ), .A2(\myexu/_1048_ ), .ZN(\myexu/_1053_ ) );
AOI21_X1 \myexu/_4056_ ( .A(\myexu/_1052_ ), .B1(\myexu/_0960_ ), .B2(\myexu/_1053_ ), .ZN(\myexu/_1054_ ) );
XNOR2_X1 \myexu/_4057_ ( .A(\myexu/_2430_ ), .B(\myexu/_2462_ ), .ZN(\myexu/_1055_ ) );
INV_X1 \myexu/_4058_ ( .A(\myexu/_1055_ ), .ZN(\myexu/_1056_ ) );
AOI21_X1 \myexu/_4059_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1054_ ), .B2(\myexu/_1056_ ), .ZN(\myexu/_1057_ ) );
OAI21_X1 \myexu/_4060_ ( .A(\myexu/_1057_ ), .B1(\myexu/_1056_ ), .B2(\myexu/_1054_ ), .ZN(\myexu/_1058_ ) );
NOR2_X1 \myexu/_4061_ ( .A1(\myexu/_0297_ ), .A2(\myexu/_2262_ ), .ZN(\myexu/_1059_ ) );
AND2_X1 \myexu/_4062_ ( .A1(\myexu/_0297_ ), .A2(\myexu/_2262_ ), .ZN(\myexu/_1060_ ) );
NOR3_X1 \myexu/_4063_ ( .A1(\myexu/_1018_ ), .A2(\myexu/_1059_ ), .A3(\myexu/_1060_ ), .ZN(\myexu/_1061_ ) );
NAND3_X1 \myexu/_4064_ ( .A1(\myexu/_0969_ ), .A2(\myexu/_1016_ ), .A3(\myexu/_1061_ ), .ZN(\myexu/_1062_ ) );
AND2_X1 \myexu/_4065_ ( .A1(\myexu/_1015_ ), .A2(\myexu/_1061_ ), .ZN(\myexu/_1063_ ) );
AND2_X1 \myexu/_4066_ ( .A1(\myexu/_1037_ ), .A2(\myexu/_1035_ ), .ZN(\myexu/_1064_ ) );
NOR3_X1 \myexu/_4067_ ( .A1(\myexu/_1063_ ), .A2(\myexu/_1060_ ), .A3(\myexu/_1064_ ), .ZN(\myexu/_1065_ ) );
AND2_X1 \myexu/_4068_ ( .A1(\myexu/_1062_ ), .A2(\myexu/_1065_ ), .ZN(\myexu/_1066_ ) );
XOR2_X1 \myexu/_4069_ ( .A(\myexu/_0298_ ), .B(\myexu/_2263_ ), .Z(\myexu/_1067_ ) );
XNOR2_X1 \myexu/_4070_ ( .A(\myexu/_1066_ ), .B(\myexu/_1067_ ), .ZN(\myexu/_1068_ ) );
AOI22_X1 \myexu/_4071_ ( .A1(\myexu/_1068_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0298_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1069_ ) );
AOI21_X1 \myexu/_4072_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1058_ ), .B2(\myexu/_1069_ ), .ZN(\myexu/_1070_ ) );
AND2_X1 \myexu/_4073_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0037_ ), .ZN(\myexu/_1071_ ) );
NOR3_X1 \myexu/_4074_ ( .A1(\myexu/_1070_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1071_ ), .ZN(\myexu/_1072_ ) );
AND3_X1 \myexu/_4075_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_2261_ ), .A3(\myexu/_2262_ ), .ZN(\myexu/_1073_ ) );
INV_X1 \myexu/_4076_ ( .A(\myexu/_2263_ ), .ZN(\myexu/_1074_ ) );
XNOR2_X1 \myexu/_4077_ ( .A(\myexu/_1073_ ), .B(\myexu/_1074_ ), .ZN(\myexu/_1075_ ) );
OAI21_X1 \myexu/_4078_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1075_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1076_ ) );
OAI221_X1 \myexu/_4079_ ( .A(\myexu/_1047_ ), .B1(\myexu/_2227_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1072_ ), .C2(\myexu/_1076_ ), .ZN(\myexu/_0221_ ) );
INV_X1 \myexu/_4080_ ( .A(\myexu/_2236_ ), .ZN(\myexu/_1077_ ) );
NOR2_X1 \myexu/_4081_ ( .A1(\myexu/_1054_ ), .A2(\myexu/_1056_ ), .ZN(\myexu/_1078_ ) );
NOR2_X1 \myexu/_4082_ ( .A1(\myexu/_2226_ ), .A2(\myexu/_2462_ ), .ZN(\myexu/_1079_ ) );
XNOR2_X1 \myexu/_4083_ ( .A(\myexu/_2431_ ), .B(\myexu/_2463_ ), .ZN(\myexu/_1080_ ) );
OR3_X1 \myexu/_4084_ ( .A1(\myexu/_1078_ ), .A2(\myexu/_1079_ ), .A3(\myexu/_1080_ ), .ZN(\myexu/_1081_ ) );
AOI21_X1 \myexu/_4085_ ( .A(\myexu/_0773_ ), .B1(\myexu/_1079_ ), .B2(\myexu/_1080_ ), .ZN(\myexu/_1082_ ) );
NAND2_X1 \myexu/_4086_ ( .A1(\myexu/_1055_ ), .A2(\myexu/_1080_ ), .ZN(\myexu/_1083_ ) );
OAI211_X2 \myexu/_4087_ ( .A(\myexu/_1081_ ), .B(\myexu/_1082_ ), .C1(\myexu/_1054_ ), .C2(\myexu/_1083_ ), .ZN(\myexu/_1084_ ) );
AND2_X1 \myexu/_4088_ ( .A1(\myexu/_0298_ ), .A2(\myexu/_2263_ ), .ZN(\myexu/_1085_ ) );
INV_X1 \myexu/_4089_ ( .A(\myexu/_1085_ ), .ZN(\myexu/_1086_ ) );
NOR2_X1 \myexu/_4090_ ( .A1(\myexu/_0298_ ), .A2(\myexu/_2263_ ), .ZN(\myexu/_1087_ ) );
OAI21_X1 \myexu/_4091_ ( .A(\myexu/_1086_ ), .B1(\myexu/_1066_ ), .B2(\myexu/_1087_ ), .ZN(\myexu/_1088_ ) );
XOR2_X1 \myexu/_4092_ ( .A(\myexu/_0299_ ), .B(\myexu/_2264_ ), .Z(\myexu/_1089_ ) );
XOR2_X1 \myexu/_4093_ ( .A(\myexu/_1088_ ), .B(\myexu/_1089_ ), .Z(\myexu/_1090_ ) );
AOI22_X1 \myexu/_4094_ ( .A1(\myexu/_1090_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0299_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1091_ ) );
AOI21_X1 \myexu/_4095_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1084_ ), .B2(\myexu/_1091_ ), .ZN(\myexu/_1092_ ) );
AND2_X1 \myexu/_4096_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0038_ ), .ZN(\myexu/_1093_ ) );
NOR3_X1 \myexu/_4097_ ( .A1(\myexu/_1092_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_1093_ ), .ZN(\myexu/_1094_ ) );
AND2_X1 \myexu/_4098_ ( .A1(\myexu/_1073_ ), .A2(\myexu/_2263_ ), .ZN(\myexu/_1095_ ) );
XNOR2_X1 \myexu/_4099_ ( .A(\myexu/_1095_ ), .B(\myexu/_2233_ ), .ZN(\myexu/_1096_ ) );
OAI21_X1 \myexu/_4100_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1096_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_1097_ ) );
OAI21_X1 \myexu/_4101_ ( .A(\myexu/_1077_ ), .B1(\myexu/_1094_ ), .B2(\myexu/_1097_ ), .ZN(\myexu/_1098_ ) );
MUX2_X1 \myexu/_4102_ ( .A(\myexu/_2398_ ), .B(\myexu/_1098_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0222_ ) );
NAND3_X1 \myexu/_4103_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_2034_ ), .A3(\myexu/_2496_ ), .ZN(\myexu/_1099_ ) );
NOR2_X1 \myexu/_4104_ ( .A1(\myexu/_0659_ ), .A2(\myexu/_2463_ ), .ZN(\myexu/_1100_ ) );
AOI21_X1 \myexu/_4105_ ( .A(\myexu/_1100_ ), .B1(\myexu/_1080_ ), .B2(\myexu/_1079_ ), .ZN(\myexu/_1101_ ) );
OAI21_X1 \myexu/_4106_ ( .A(\myexu/_1101_ ), .B1(\myexu/_1054_ ), .B2(\myexu/_1083_ ), .ZN(\myexu/_1102_ ) );
XNOR2_X1 \myexu/_4107_ ( .A(\myexu/_2432_ ), .B(\myexu/_2464_ ), .ZN(\myexu/_1103_ ) );
AND2_X1 \myexu/_4108_ ( .A1(\myexu/_1102_ ), .A2(\myexu/_1103_ ), .ZN(\myexu/_1104_ ) );
OAI21_X1 \myexu/_4109_ ( .A(\myexu/_0834_ ), .B1(\myexu/_1102_ ), .B2(\myexu/_1103_ ), .ZN(\myexu/_1105_ ) );
OR2_X1 \myexu/_4110_ ( .A1(\myexu/_1104_ ), .A2(\myexu/_1105_ ), .ZN(\myexu/_1106_ ) );
AND2_X1 \myexu/_4111_ ( .A1(\myexu/_0299_ ), .A2(\myexu/_2264_ ), .ZN(\myexu/_1107_ ) );
AOI21_X1 \myexu/_4112_ ( .A(\myexu/_1107_ ), .B1(\myexu/_1088_ ), .B2(\myexu/_1089_ ), .ZN(\myexu/_1108_ ) );
XNOR2_X1 \myexu/_4113_ ( .A(\myexu/_0300_ ), .B(\myexu/_2265_ ), .ZN(\myexu/_1109_ ) );
XOR2_X1 \myexu/_4114_ ( .A(\myexu/_1108_ ), .B(\myexu/_1109_ ), .Z(\myexu/_1110_ ) );
AOI22_X1 \myexu/_4115_ ( .A1(\myexu/_1110_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0300_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1111_ ) );
AOI21_X1 \myexu/_4116_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1106_ ), .B2(\myexu/_1111_ ), .ZN(\myexu/_1112_ ) );
AND2_X1 \myexu/_4117_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0039_ ), .ZN(\myexu/_1113_ ) );
NOR3_X1 \myexu/_4118_ ( .A1(\myexu/_1112_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_1113_ ), .ZN(\myexu/_1114_ ) );
AND2_X1 \myexu/_4119_ ( .A1(\myexu/_2263_ ), .A2(\myexu/_2264_ ), .ZN(\myexu/_1115_ ) );
AND3_X1 \myexu/_4120_ ( .A1(\myexu/_1115_ ), .A2(\myexu/_2261_ ), .A3(\myexu/_2262_ ), .ZN(\myexu/_1116_ ) );
AND2_X4 \myexu/_4121_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_1116_ ), .ZN(\myexu/_1117_ ) );
INV_X1 \myexu/_4122_ ( .A(\myexu/_2265_ ), .ZN(\myexu/_1118_ ) );
XNOR2_X1 \myexu/_4123_ ( .A(\myexu/_1117_ ), .B(\myexu/_1118_ ), .ZN(\myexu/_1119_ ) );
OAI21_X1 \myexu/_4124_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1119_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_1120_ ) );
OAI21_X1 \myexu/_4125_ ( .A(\myexu/_1099_ ), .B1(\myexu/_1114_ ), .B2(\myexu/_1120_ ), .ZN(\myexu/_1121_ ) );
MUX2_X1 \myexu/_4126_ ( .A(\myexu/_2399_ ), .B(\myexu/_1121_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0223_ ) );
OAI21_X1 \myexu/_4127_ ( .A(\myexu/_2400_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1122_ ) );
NOR2_X1 \myexu/_4128_ ( .A1(\myexu/_0655_ ), .A2(\myexu/_2464_ ), .ZN(\myexu/_1123_ ) );
XNOR2_X1 \myexu/_4129_ ( .A(\myexu/_2433_ ), .B(\myexu/_2465_ ), .ZN(\myexu/_1124_ ) );
OR3_X1 \myexu/_4130_ ( .A1(\myexu/_1104_ ), .A2(\myexu/_1123_ ), .A3(\myexu/_1124_ ), .ZN(\myexu/_1125_ ) );
OAI21_X1 \myexu/_4131_ ( .A(\myexu/_1124_ ), .B1(\myexu/_1104_ ), .B2(\myexu/_1123_ ), .ZN(\myexu/_1126_ ) );
NAND3_X1 \myexu/_4132_ ( .A1(\myexu/_1125_ ), .A2(\myexu/_0834_ ), .A3(\myexu/_1126_ ), .ZN(\myexu/_1127_ ) );
NOR2_X1 \myexu/_4133_ ( .A1(\myexu/_1108_ ), .A2(\myexu/_1109_ ), .ZN(\myexu/_1128_ ) );
AND2_X1 \myexu/_4134_ ( .A1(\myexu/_0300_ ), .A2(\myexu/_2265_ ), .ZN(\myexu/_1129_ ) );
NOR2_X1 \myexu/_4135_ ( .A1(\myexu/_1128_ ), .A2(\myexu/_1129_ ), .ZN(\myexu/_1130_ ) );
XOR2_X1 \myexu/_4136_ ( .A(\myexu/_0301_ ), .B(\myexu/_2266_ ), .Z(\myexu/_1131_ ) );
XNOR2_X1 \myexu/_4137_ ( .A(\myexu/_1130_ ), .B(\myexu/_1131_ ), .ZN(\myexu/_1132_ ) );
AOI22_X1 \myexu/_4138_ ( .A1(\myexu/_1132_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0301_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1133_ ) );
AOI21_X1 \myexu/_4139_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1127_ ), .B2(\myexu/_1133_ ), .ZN(\myexu/_1134_ ) );
AND2_X1 \myexu/_4140_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0040_ ), .ZN(\myexu/_1135_ ) );
NOR3_X1 \myexu/_4141_ ( .A1(\myexu/_1134_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1135_ ), .ZN(\myexu/_1136_ ) );
AND2_X1 \myexu/_4142_ ( .A1(\myexu/_1117_ ), .A2(\myexu/_2265_ ), .ZN(\myexu/_1137_ ) );
XNOR2_X1 \myexu/_4143_ ( .A(\myexu/_1137_ ), .B(\myexu/_2256_ ), .ZN(\myexu/_1138_ ) );
OAI21_X1 \myexu/_4144_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1138_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1139_ ) );
OAI221_X1 \myexu/_4145_ ( .A(\myexu/_1122_ ), .B1(\myexu/_2251_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1136_ ), .C2(\myexu/_1139_ ), .ZN(\myexu/_0224_ ) );
NAND3_X1 \myexu/_4146_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_1963_ ), .A3(\myexu/_2498_ ), .ZN(\myexu/_1140_ ) );
NAND2_X1 \myexu/_4147_ ( .A1(\myexu/_1103_ ), .A2(\myexu/_1124_ ), .ZN(\myexu/_1141_ ) );
NOR2_X1 \myexu/_4148_ ( .A1(\myexu/_1083_ ), .A2(\myexu/_1141_ ), .ZN(\myexu/_1142_ ) );
AND3_X4 \myexu/_4149_ ( .A1(\myexu/_0960_ ), .A2(\myexu/_1053_ ), .A3(\myexu/_1142_ ), .ZN(\myexu/_1143_ ) );
AND2_X1 \myexu/_4150_ ( .A1(\myexu/_1052_ ), .A2(\myexu/_1142_ ), .ZN(\myexu/_1144_ ) );
AND2_X1 \myexu/_4151_ ( .A1(\myexu/_2255_ ), .A2(\myexu/_2433_ ), .ZN(\myexu/_1145_ ) );
NOR2_X1 \myexu/_4152_ ( .A1(\myexu/_1101_ ), .A2(\myexu/_1141_ ), .ZN(\myexu/_1146_ ) );
AND2_X1 \myexu/_4153_ ( .A1(\myexu/_1124_ ), .A2(\myexu/_1123_ ), .ZN(\myexu/_1147_ ) );
NOR4_X1 \myexu/_4154_ ( .A1(\myexu/_1144_ ), .A2(\myexu/_1145_ ), .A3(\myexu/_1146_ ), .A4(\myexu/_1147_ ), .ZN(\myexu/_1148_ ) );
INV_X1 \myexu/_4155_ ( .A(\myexu/_1148_ ), .ZN(\myexu/_1149_ ) );
NOR2_X1 \myexu/_4156_ ( .A1(\myexu/_1143_ ), .A2(\myexu/_1149_ ), .ZN(\myexu/_1150_ ) );
INV_X1 \myexu/_4157_ ( .A(\myexu/_1150_ ), .ZN(\myexu/_1151_ ) );
XNOR2_X1 \myexu/_4158_ ( .A(\myexu/_2434_ ), .B(\myexu/_2466_ ), .ZN(\myexu/_1152_ ) );
AOI21_X1 \myexu/_4159_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1151_ ), .B2(\myexu/_1152_ ), .ZN(\myexu/_1153_ ) );
OAI21_X1 \myexu/_4160_ ( .A(\myexu/_1153_ ), .B1(\myexu/_1151_ ), .B2(\myexu/_1152_ ), .ZN(\myexu/_1154_ ) );
INV_X1 \myexu/_4161_ ( .A(\myexu/_1131_ ), .ZN(\myexu/_1155_ ) );
NOR4_X1 \myexu/_4162_ ( .A1(\myexu/_1155_ ), .A2(\myexu/_1087_ ), .A3(\myexu/_1085_ ), .A4(\myexu/_1109_ ), .ZN(\myexu/_1156_ ) );
NAND2_X1 \myexu/_4163_ ( .A1(\myexu/_1156_ ), .A2(\myexu/_1089_ ), .ZN(\myexu/_1157_ ) );
OR2_X1 \myexu/_4164_ ( .A1(\myexu/_1062_ ), .A2(\myexu/_1157_ ), .ZN(\myexu/_1158_ ) );
AND2_X1 \myexu/_4165_ ( .A1(\myexu/_1131_ ), .A2(\myexu/_1129_ ), .ZN(\myexu/_1159_ ) );
AOI21_X1 \myexu/_4166_ ( .A(\myexu/_1107_ ), .B1(\myexu/_1089_ ), .B2(\myexu/_1085_ ), .ZN(\myexu/_1160_ ) );
OR3_X1 \myexu/_4167_ ( .A1(\myexu/_1160_ ), .A2(\myexu/_1109_ ), .A3(\myexu/_1155_ ), .ZN(\myexu/_1161_ ) );
OAI21_X1 \myexu/_4168_ ( .A(\myexu/_1161_ ), .B1(\myexu/_1065_ ), .B2(\myexu/_1157_ ), .ZN(\myexu/_1162_ ) );
AOI211_X4 \myexu/_4169_ ( .A(\myexu/_1159_ ), .B(\myexu/_1162_ ), .C1(\myexu/_0301_ ), .C2(\myexu/_2266_ ), .ZN(\myexu/_1163_ ) );
NAND2_X2 \myexu/_4170_ ( .A1(\myexu/_1158_ ), .A2(\myexu/_1163_ ), .ZN(\myexu/_1164_ ) );
XOR2_X1 \myexu/_4171_ ( .A(\myexu/_0302_ ), .B(\myexu/_2267_ ), .Z(\myexu/_1165_ ) );
XOR2_X1 \myexu/_4172_ ( .A(\myexu/_1164_ ), .B(\myexu/_1165_ ), .Z(\myexu/_1166_ ) );
AOI22_X1 \myexu/_4173_ ( .A1(\myexu/_1166_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0302_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1167_ ) );
AOI21_X1 \myexu/_4174_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1154_ ), .B2(\myexu/_1167_ ), .ZN(\myexu/_1168_ ) );
AND2_X1 \myexu/_4175_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0041_ ), .ZN(\myexu/_1169_ ) );
NOR3_X1 \myexu/_4176_ ( .A1(\myexu/_1168_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_1169_ ), .ZN(\myexu/_1170_ ) );
AND2_X1 \myexu/_4177_ ( .A1(\myexu/_2265_ ), .A2(\myexu/_2266_ ), .ZN(\myexu/_1171_ ) );
NAND3_X1 \myexu/_4178_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_1116_ ), .A3(\myexu/_1171_ ), .ZN(\myexu/_1172_ ) );
XNOR2_X1 \myexu/_4179_ ( .A(\myexu/_1172_ ), .B(\myexu/_2267_ ), .ZN(\myexu/_1173_ ) );
OAI21_X1 \myexu/_4180_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1173_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_1174_ ) );
OAI21_X1 \myexu/_4181_ ( .A(\myexu/_1140_ ), .B1(\myexu/_1170_ ), .B2(\myexu/_1174_ ), .ZN(\myexu/_1175_ ) );
MUX2_X1 \myexu/_4182_ ( .A(\myexu/_2401_ ), .B(\myexu/_1175_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0225_ ) );
NOR2_X1 \myexu/_4183_ ( .A1(\myexu/_0723_ ), .A2(\myexu/_2466_ ), .ZN(\myexu/_1176_ ) );
AOI21_X1 \myexu/_4184_ ( .A(\myexu/_1176_ ), .B1(\myexu/_1151_ ), .B2(\myexu/_1152_ ), .ZN(\myexu/_1177_ ) );
XNOR2_X1 \myexu/_4185_ ( .A(\myexu/_2435_ ), .B(\myexu/_2467_ ), .ZN(\myexu/_1178_ ) );
XNOR2_X1 \myexu/_4186_ ( .A(\myexu/_1177_ ), .B(\myexu/_1178_ ), .ZN(\myexu/_1179_ ) );
AND3_X1 \myexu/_4187_ ( .A1(\myexu/_1179_ ), .A2(\myexu/_0770_ ), .A3(\myexu/_0763_ ), .ZN(\myexu/_1180_ ) );
AND3_X1 \myexu/_4188_ ( .A1(\myexu/_0776_ ), .A2(\myexu/_0777_ ), .A3(\myexu/_0303_ ), .ZN(\myexu/_1181_ ) );
OR2_X1 \myexu/_4189_ ( .A1(\myexu/_1180_ ), .A2(\myexu/_1181_ ), .ZN(\myexu/_1182_ ) );
NAND2_X1 \myexu/_4190_ ( .A1(\myexu/_1164_ ), .A2(\myexu/_1165_ ), .ZN(\myexu/_1183_ ) );
AND2_X1 \myexu/_4191_ ( .A1(\myexu/_0302_ ), .A2(\myexu/_2267_ ), .ZN(\myexu/_1184_ ) );
INV_X1 \myexu/_4192_ ( .A(\myexu/_1184_ ), .ZN(\myexu/_1185_ ) );
AND2_X1 \myexu/_4193_ ( .A1(\myexu/_1183_ ), .A2(\myexu/_1185_ ), .ZN(\myexu/_1186_ ) );
AND2_X1 \myexu/_4194_ ( .A1(\myexu/_0303_ ), .A2(\myexu/_2268_ ), .ZN(\myexu/_1187_ ) );
NOR2_X1 \myexu/_4195_ ( .A1(\myexu/_0303_ ), .A2(\myexu/_2268_ ), .ZN(\myexu/_1188_ ) );
NOR2_X1 \myexu/_4196_ ( .A1(\myexu/_1187_ ), .A2(\myexu/_1188_ ), .ZN(\myexu/_1189_ ) );
XNOR2_X1 \myexu/_4197_ ( .A(\myexu/_1186_ ), .B(\myexu/_1189_ ), .ZN(\myexu/_1190_ ) );
AND2_X1 \myexu/_4198_ ( .A1(\myexu/_1190_ ), .A2(\myexu/_0780_ ), .ZN(\myexu/_1191_ ) );
OAI21_X1 \myexu/_4199_ ( .A(\myexu/_0800_ ), .B1(\myexu/_1182_ ), .B2(\myexu/_1191_ ), .ZN(\myexu/_1192_ ) );
AOI21_X1 \myexu/_4200_ ( .A(\myexu/_0785_ ), .B1(\myexu/_0791_ ), .B2(\myexu/_0042_ ), .ZN(\myexu/_1193_ ) );
INV_X1 \myexu/_4201_ ( .A(\myexu/_2267_ ), .ZN(\myexu/_1194_ ) );
NOR2_X1 \myexu/_4202_ ( .A1(\myexu/_1172_ ), .A2(\myexu/_1194_ ), .ZN(\myexu/_1195_ ) );
XNOR2_X1 \myexu/_4203_ ( .A(\myexu/_1195_ ), .B(\myexu/_2268_ ), .ZN(\myexu/_1196_ ) );
AOI22_X1 \myexu/_4204_ ( .A1(\myexu/_1192_ ), .A2(\myexu/_1193_ ), .B1(\myexu/_0786_ ), .B2(\myexu/_1196_ ), .ZN(\myexu/_1197_ ) );
MUX2_X1 \myexu/_4205_ ( .A(\myexu/_2499_ ), .B(\myexu/_1197_ ), .S(\myexu/_2131_ ), .Z(\myexu/_1198_ ) );
MUX2_X1 \myexu/_4206_ ( .A(\myexu/_2402_ ), .B(\myexu/_1198_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0226_ ) );
OAI21_X1 \myexu/_4207_ ( .A(\myexu/_2403_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1199_ ) );
NAND4_X1 \myexu/_4208_ ( .A1(\myexu/_2049_ ), .A2(\myexu/_1972_ ), .A3(\myexu/_2500_ ), .A4(\myexu/_2003_ ), .ZN(\myexu/_1200_ ) );
AND2_X1 \myexu/_4209_ ( .A1(\myexu/_1178_ ), .A2(\myexu/_1176_ ), .ZN(\myexu/_1201_ ) );
INV_X1 \myexu/_4210_ ( .A(\myexu/_1201_ ), .ZN(\myexu/_1202_ ) );
OAI21_X1 \myexu/_4211_ ( .A(\myexu/_1202_ ), .B1(\myexu/_0333_ ), .B2(\myexu/_2467_ ), .ZN(\myexu/_1203_ ) );
AND2_X1 \myexu/_4212_ ( .A1(\myexu/_1152_ ), .A2(\myexu/_1178_ ), .ZN(\myexu/_1204_ ) );
AOI21_X1 \myexu/_4213_ ( .A(\myexu/_1203_ ), .B1(\myexu/_1151_ ), .B2(\myexu/_1204_ ), .ZN(\myexu/_1205_ ) );
XNOR2_X1 \myexu/_4214_ ( .A(\myexu/_2436_ ), .B(\myexu/_2468_ ), .ZN(\myexu/_1206_ ) );
INV_X1 \myexu/_4215_ ( .A(\myexu/_1206_ ), .ZN(\myexu/_1207_ ) );
AOI21_X1 \myexu/_4216_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1205_ ), .B2(\myexu/_1207_ ), .ZN(\myexu/_1208_ ) );
OAI21_X1 \myexu/_4217_ ( .A(\myexu/_1208_ ), .B1(\myexu/_1205_ ), .B2(\myexu/_1207_ ), .ZN(\myexu/_1209_ ) );
AOI21_X1 \myexu/_4218_ ( .A(\myexu/_1187_ ), .B1(\myexu/_1189_ ), .B2(\myexu/_1184_ ), .ZN(\myexu/_1210_ ) );
INV_X1 \myexu/_4219_ ( .A(\myexu/_1210_ ), .ZN(\myexu/_1211_ ) );
AND2_X1 \myexu/_4220_ ( .A1(\myexu/_1165_ ), .A2(\myexu/_1189_ ), .ZN(\myexu/_1212_ ) );
AOI21_X1 \myexu/_4221_ ( .A(\myexu/_1211_ ), .B1(\myexu/_1164_ ), .B2(\myexu/_1212_ ), .ZN(\myexu/_1213_ ) );
XOR2_X1 \myexu/_4222_ ( .A(\myexu/_0304_ ), .B(\myexu/_2269_ ), .Z(\myexu/_1214_ ) );
XNOR2_X1 \myexu/_4223_ ( .A(\myexu/_1213_ ), .B(\myexu/_1214_ ), .ZN(\myexu/_1215_ ) );
AOI22_X1 \myexu/_4224_ ( .A1(\myexu/_1215_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0304_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1216_ ) );
AOI21_X1 \myexu/_4225_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1209_ ), .B2(\myexu/_1216_ ), .ZN(\myexu/_1217_ ) );
AND2_X1 \myexu/_4226_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0043_ ), .ZN(\myexu/_1218_ ) );
NOR3_X1 \myexu/_4227_ ( .A1(\myexu/_1217_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1218_ ), .ZN(\myexu/_1219_ ) );
AND4_X1 \myexu/_4228_ ( .A1(\myexu/_2267_ ), .A2(\myexu/_1116_ ), .A3(\myexu/_2268_ ), .A4(\myexu/_1171_ ), .ZN(\myexu/_1220_ ) );
NAND2_X1 \myexu/_4229_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_1220_ ), .ZN(\myexu/_1221_ ) );
XNOR2_X1 \myexu/_4230_ ( .A(\myexu/_1221_ ), .B(\myexu/_2269_ ), .ZN(\myexu/_1222_ ) );
OAI21_X1 \myexu/_4231_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1222_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1223_ ) );
OAI211_X2 \myexu/_4232_ ( .A(\myexu/_1199_ ), .B(\myexu/_1200_ ), .C1(\myexu/_1219_ ), .C2(\myexu/_1223_ ), .ZN(\myexu/_0227_ ) );
OAI21_X1 \myexu/_4233_ ( .A(\myexu/_2404_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1224_ ) );
NOR2_X1 \myexu/_4234_ ( .A1(\myexu/_0342_ ), .A2(\myexu/_2468_ ), .ZN(\myexu/_1225_ ) );
INV_X1 \myexu/_4235_ ( .A(\myexu/_1225_ ), .ZN(\myexu/_1226_ ) );
OAI21_X1 \myexu/_4236_ ( .A(\myexu/_1226_ ), .B1(\myexu/_1205_ ), .B2(\myexu/_1207_ ), .ZN(\myexu/_1227_ ) );
XNOR2_X1 \myexu/_4237_ ( .A(\myexu/_2437_ ), .B(\myexu/_2469_ ), .ZN(\myexu/_1228_ ) );
AOI21_X1 \myexu/_4238_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1227_ ), .B2(\myexu/_1228_ ), .ZN(\myexu/_1229_ ) );
OAI21_X1 \myexu/_4239_ ( .A(\myexu/_1229_ ), .B1(\myexu/_1227_ ), .B2(\myexu/_1228_ ), .ZN(\myexu/_1230_ ) );
NOR2_X1 \myexu/_4240_ ( .A1(\myexu/_0304_ ), .A2(\myexu/_2269_ ), .ZN(\myexu/_1231_ ) );
AND2_X1 \myexu/_4241_ ( .A1(\myexu/_0304_ ), .A2(\myexu/_2269_ ), .ZN(\myexu/_1232_ ) );
NOR3_X1 \myexu/_4242_ ( .A1(\myexu/_1213_ ), .A2(\myexu/_1231_ ), .A3(\myexu/_1232_ ), .ZN(\myexu/_1233_ ) );
NOR2_X1 \myexu/_4243_ ( .A1(\myexu/_1233_ ), .A2(\myexu/_1232_ ), .ZN(\myexu/_1234_ ) );
XOR2_X1 \myexu/_4244_ ( .A(\myexu/_0305_ ), .B(\myexu/_2270_ ), .Z(\myexu/_1235_ ) );
XNOR2_X1 \myexu/_4245_ ( .A(\myexu/_1234_ ), .B(\myexu/_1235_ ), .ZN(\myexu/_1236_ ) );
AOI22_X1 \myexu/_4246_ ( .A1(\myexu/_1236_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0305_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1237_ ) );
AOI21_X1 \myexu/_4247_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1230_ ), .B2(\myexu/_1237_ ), .ZN(\myexu/_1238_ ) );
AND2_X1 \myexu/_4248_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0044_ ), .ZN(\myexu/_1239_ ) );
NOR3_X1 \myexu/_4249_ ( .A1(\myexu/_1238_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1239_ ), .ZN(\myexu/_1240_ ) );
NAND3_X1 \myexu/_4250_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_2269_ ), .A3(\myexu/_1220_ ), .ZN(\myexu/_1241_ ) );
XNOR2_X1 \myexu/_4251_ ( .A(\myexu/_1241_ ), .B(\myexu/_2270_ ), .ZN(\myexu/_1242_ ) );
OAI21_X1 \myexu/_4252_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1242_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1243_ ) );
OAI221_X1 \myexu/_4253_ ( .A(\myexu/_1224_ ), .B1(\myexu/_0349_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1240_ ), .C2(\myexu/_1243_ ), .ZN(\myexu/_0228_ ) );
AND2_X1 \myexu/_4254_ ( .A1(\myexu/_1206_ ), .A2(\myexu/_1228_ ), .ZN(\myexu/_1244_ ) );
AND2_X1 \myexu/_4255_ ( .A1(\myexu/_1203_ ), .A2(\myexu/_1244_ ), .ZN(\myexu/_1245_ ) );
NOR2_X1 \myexu/_4256_ ( .A1(\myexu/_0348_ ), .A2(\myexu/_2469_ ), .ZN(\myexu/_1246_ ) );
AND2_X1 \myexu/_4257_ ( .A1(\myexu/_1228_ ), .A2(\myexu/_1225_ ), .ZN(\myexu/_1247_ ) );
NOR3_X1 \myexu/_4258_ ( .A1(\myexu/_1245_ ), .A2(\myexu/_1246_ ), .A3(\myexu/_1247_ ), .ZN(\myexu/_1248_ ) );
NAND2_X1 \myexu/_4259_ ( .A1(\myexu/_1204_ ), .A2(\myexu/_1244_ ), .ZN(\myexu/_1249_ ) );
OAI21_X1 \myexu/_4260_ ( .A(\myexu/_1248_ ), .B1(\myexu/_1150_ ), .B2(\myexu/_1249_ ), .ZN(\myexu/_1250_ ) );
XNOR2_X1 \myexu/_4261_ ( .A(\myexu/_2439_ ), .B(\myexu/_2471_ ), .ZN(\myexu/_1251_ ) );
AOI21_X1 \myexu/_4262_ ( .A(\myexu/_0773_ ), .B1(\myexu/_1250_ ), .B2(\myexu/_1251_ ), .ZN(\myexu/_1252_ ) );
OAI21_X1 \myexu/_4263_ ( .A(\myexu/_1252_ ), .B1(\myexu/_1251_ ), .B2(\myexu/_1250_ ), .ZN(\myexu/_1253_ ) );
AND2_X1 \myexu/_4264_ ( .A1(\myexu/_1214_ ), .A2(\myexu/_1235_ ), .ZN(\myexu/_1254_ ) );
NAND3_X1 \myexu/_4265_ ( .A1(\myexu/_1164_ ), .A2(\myexu/_1212_ ), .A3(\myexu/_1254_ ), .ZN(\myexu/_1255_ ) );
AND2_X1 \myexu/_4266_ ( .A1(\myexu/_1211_ ), .A2(\myexu/_1254_ ), .ZN(\myexu/_1256_ ) );
AND2_X1 \myexu/_4267_ ( .A1(\myexu/_0305_ ), .A2(\myexu/_2270_ ), .ZN(\myexu/_1257_ ) );
AND2_X1 \myexu/_4268_ ( .A1(\myexu/_1235_ ), .A2(\myexu/_1232_ ), .ZN(\myexu/_1258_ ) );
NOR3_X1 \myexu/_4269_ ( .A1(\myexu/_1256_ ), .A2(\myexu/_1257_ ), .A3(\myexu/_1258_ ), .ZN(\myexu/_1259_ ) );
AND2_X1 \myexu/_4270_ ( .A1(\myexu/_1255_ ), .A2(\myexu/_1259_ ), .ZN(\myexu/_1260_ ) );
XOR2_X1 \myexu/_4271_ ( .A(\myexu/_0307_ ), .B(\myexu/_2272_ ), .Z(\myexu/_1261_ ) );
XNOR2_X1 \myexu/_4272_ ( .A(\myexu/_1260_ ), .B(\myexu/_1261_ ), .ZN(\myexu/_1262_ ) );
AOI22_X1 \myexu/_4273_ ( .A1(\myexu/_1262_ ), .A2(\myexu/_0780_ ), .B1(\myexu/_0307_ ), .B2(\myexu/_0778_ ), .ZN(\myexu/_1263_ ) );
AOI21_X1 \myexu/_4274_ ( .A(\myexu/_0639_ ), .B1(\myexu/_1253_ ), .B2(\myexu/_1263_ ), .ZN(\myexu/_1264_ ) );
AND2_X1 \myexu/_4275_ ( .A1(\myexu/_0791_ ), .A2(\myexu/_0046_ ), .ZN(\myexu/_1265_ ) );
NOR3_X1 \myexu/_4276_ ( .A1(\myexu/_1264_ ), .A2(\myexu/_0785_ ), .A3(\myexu/_1265_ ), .ZN(\myexu/_1266_ ) );
BUF_X4 \myexu/_4277_ ( .A(\myexu/_0785_ ), .Z(\myexu/_1267_ ) );
NAND2_X1 \myexu/_4278_ ( .A1(\myexu/_2269_ ), .A2(\myexu/_2270_ ), .ZN(\myexu/_1268_ ) );
NOR2_X1 \myexu/_4279_ ( .A1(\myexu/_1221_ ), .A2(\myexu/_1268_ ), .ZN(\myexu/_1269_ ) );
XNOR2_X1 \myexu/_4280_ ( .A(\myexu/_1269_ ), .B(\myexu/_2272_ ), .ZN(\myexu/_1270_ ) );
AOI21_X1 \myexu/_4281_ ( .A(\myexu/_1266_ ), .B1(\myexu/_1267_ ), .B2(\myexu/_1270_ ), .ZN(\myexu/_1271_ ) );
MUX2_X1 \myexu/_4282_ ( .A(\myexu/_2503_ ), .B(\myexu/_1271_ ), .S(\myexu/_2131_ ), .Z(\myexu/_1272_ ) );
MUX2_X1 \myexu/_4283_ ( .A(\myexu/_2406_ ), .B(\myexu/_1272_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0229_ ) );
INV_X1 \myexu/_4284_ ( .A(\myexu/_2272_ ), .ZN(\myexu/_1273_ ) );
NOR3_X1 \myexu/_4285_ ( .A1(\myexu/_1221_ ), .A2(\myexu/_1273_ ), .A3(\myexu/_1268_ ), .ZN(\myexu/_1274_ ) );
XNOR2_X1 \myexu/_4286_ ( .A(\myexu/_1274_ ), .B(\myexu/_0364_ ), .ZN(\myexu/_1275_ ) );
NOR2_X1 \myexu/_4287_ ( .A1(\myexu/_1275_ ), .A2(\myexu/_0795_ ), .ZN(\myexu/_1276_ ) );
AND2_X1 \myexu/_4288_ ( .A1(\myexu/_1250_ ), .A2(\myexu/_1251_ ), .ZN(\myexu/_1277_ ) );
NOR2_X1 \myexu/_4289_ ( .A1(\myexu/_0714_ ), .A2(\myexu/_2471_ ), .ZN(\myexu/_1278_ ) );
XNOR2_X1 \myexu/_4290_ ( .A(\myexu/_2440_ ), .B(\myexu/_2472_ ), .ZN(\myexu/_1279_ ) );
NOR3_X1 \myexu/_4291_ ( .A1(\myexu/_1277_ ), .A2(\myexu/_1278_ ), .A3(\myexu/_1279_ ), .ZN(\myexu/_1280_ ) );
AND2_X1 \myexu/_4292_ ( .A1(\myexu/_1279_ ), .A2(\myexu/_1278_ ), .ZN(\myexu/_1281_ ) );
OR3_X1 \myexu/_4293_ ( .A1(\myexu/_1280_ ), .A2(\myexu/_0773_ ), .A3(\myexu/_1281_ ), .ZN(\myexu/_1282_ ) );
AOI21_X1 \myexu/_4294_ ( .A(\myexu/_1282_ ), .B1(\myexu/_1277_ ), .B2(\myexu/_1279_ ), .ZN(\myexu/_1283_ ) );
INV_X1 \myexu/_4295_ ( .A(\myexu/_1261_ ), .ZN(\myexu/_1284_ ) );
AOI21_X1 \myexu/_4296_ ( .A(\myexu/_1284_ ), .B1(\myexu/_1255_ ), .B2(\myexu/_1259_ ), .ZN(\myexu/_1285_ ) );
INV_X1 \myexu/_4297_ ( .A(\myexu/_1285_ ), .ZN(\myexu/_1286_ ) );
NAND2_X1 \myexu/_4298_ ( .A1(\myexu/_0307_ ), .A2(\myexu/_2272_ ), .ZN(\myexu/_1287_ ) );
NAND2_X1 \myexu/_4299_ ( .A1(\myexu/_1286_ ), .A2(\myexu/_1287_ ), .ZN(\myexu/_1288_ ) );
XOR2_X1 \myexu/_4300_ ( .A(\myexu/_0308_ ), .B(\myexu/_2273_ ), .Z(\myexu/_1289_ ) );
INV_X1 \myexu/_4301_ ( .A(\myexu/_1289_ ), .ZN(\myexu/_1290_ ) );
XNOR2_X1 \myexu/_4302_ ( .A(\myexu/_1288_ ), .B(\myexu/_1290_ ), .ZN(\myexu/_1291_ ) );
NAND2_X1 \myexu/_4303_ ( .A1(\myexu/_1291_ ), .A2(\myexu/_0780_ ), .ZN(\myexu/_1292_ ) );
INV_X1 \myexu/_4304_ ( .A(\myexu/_0308_ ), .ZN(\myexu/_1293_ ) );
OAI21_X1 \myexu/_4305_ ( .A(\myexu/_1292_ ), .B1(\myexu/_1293_ ), .B2(\myexu/_0806_ ), .ZN(\myexu/_1294_ ) );
OAI21_X1 \myexu/_4306_ ( .A(\myexu/_0800_ ), .B1(\myexu/_1283_ ), .B2(\myexu/_1294_ ), .ZN(\myexu/_1295_ ) );
AOI21_X1 \myexu/_4307_ ( .A(\myexu/_0786_ ), .B1(\myexu/_0885_ ), .B2(\myexu/_0047_ ), .ZN(\myexu/_1296_ ) );
AOI21_X1 \myexu/_4308_ ( .A(\myexu/_1276_ ), .B1(\myexu/_1295_ ), .B2(\myexu/_1296_ ), .ZN(\myexu/_1297_ ) );
MUX2_X1 \myexu/_4309_ ( .A(\myexu/_2504_ ), .B(\myexu/_1297_ ), .S(\myexu/_2131_ ), .Z(\myexu/_1298_ ) );
MUX2_X1 \myexu/_4310_ ( .A(\myexu/_2407_ ), .B(\myexu/_1298_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0230_ ) );
OAI21_X1 \myexu/_4311_ ( .A(\myexu/_2408_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1299_ ) );
INV_X1 \myexu/_4312_ ( .A(\myexu/_2505_ ), .ZN(\myexu/_1300_ ) );
AOI21_X1 \myexu/_4313_ ( .A(\myexu/_1281_ ), .B1(\myexu/_2440_ ), .B2(\myexu/_0363_ ), .ZN(\myexu/_1301_ ) );
INV_X1 \myexu/_4314_ ( .A(\myexu/_1301_ ), .ZN(\myexu/_1302_ ) );
AND2_X1 \myexu/_4315_ ( .A1(\myexu/_1251_ ), .A2(\myexu/_1279_ ), .ZN(\myexu/_1303_ ) );
AOI21_X1 \myexu/_4316_ ( .A(\myexu/_1302_ ), .B1(\myexu/_1250_ ), .B2(\myexu/_1303_ ), .ZN(\myexu/_1304_ ) );
XNOR2_X1 \myexu/_4317_ ( .A(\myexu/_2441_ ), .B(\myexu/_2473_ ), .ZN(\myexu/_1305_ ) );
INV_X1 \myexu/_4318_ ( .A(\myexu/_1305_ ), .ZN(\myexu/_1306_ ) );
AOI21_X1 \myexu/_4319_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1304_ ), .B2(\myexu/_1306_ ), .ZN(\myexu/_1307_ ) );
OAI21_X1 \myexu/_4320_ ( .A(\myexu/_1307_ ), .B1(\myexu/_1304_ ), .B2(\myexu/_1306_ ), .ZN(\myexu/_1308_ ) );
NOR2_X1 \myexu/_4321_ ( .A1(\myexu/_0308_ ), .A2(\myexu/_2273_ ), .ZN(\myexu/_1309_ ) );
INV_X1 \myexu/_4322_ ( .A(\myexu/_1309_ ), .ZN(\myexu/_1310_ ) );
OAI21_X1 \myexu/_4323_ ( .A(\myexu/_1287_ ), .B1(\myexu/_1293_ ), .B2(\myexu/_0364_ ), .ZN(\myexu/_1311_ ) );
OAI21_X1 \myexu/_4324_ ( .A(\myexu/_1310_ ), .B1(\myexu/_1285_ ), .B2(\myexu/_1311_ ), .ZN(\myexu/_1312_ ) );
XOR2_X1 \myexu/_4325_ ( .A(\myexu/_0309_ ), .B(\myexu/_2274_ ), .Z(\myexu/_1313_ ) );
XNOR2_X1 \myexu/_4326_ ( .A(\myexu/_1312_ ), .B(\myexu/_1313_ ), .ZN(\myexu/_1314_ ) );
AOI22_X1 \myexu/_4327_ ( .A1(\myexu/_1314_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0309_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1315_ ) );
AOI21_X1 \myexu/_4328_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1308_ ), .B2(\myexu/_1315_ ), .ZN(\myexu/_1316_ ) );
AND2_X1 \myexu/_4329_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0048_ ), .ZN(\myexu/_1317_ ) );
NOR3_X1 \myexu/_4330_ ( .A1(\myexu/_1316_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1317_ ), .ZN(\myexu/_1318_ ) );
AND2_X1 \myexu/_4331_ ( .A1(\myexu/_1024_ ), .A2(\myexu/_1220_ ), .ZN(\myexu/_1319_ ) );
NOR3_X1 \myexu/_4332_ ( .A1(\myexu/_1268_ ), .A2(\myexu/_1273_ ), .A3(\myexu/_0364_ ), .ZN(\myexu/_1320_ ) );
NAND2_X1 \myexu/_4333_ ( .A1(\myexu/_1319_ ), .A2(\myexu/_1320_ ), .ZN(\myexu/_1321_ ) );
XNOR2_X1 \myexu/_4334_ ( .A(\myexu/_1321_ ), .B(\myexu/_2274_ ), .ZN(\myexu/_1322_ ) );
OAI21_X1 \myexu/_4335_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1322_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1323_ ) );
OAI221_X1 \myexu/_4336_ ( .A(\myexu/_1299_ ), .B1(\myexu/_1300_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1318_ ), .C2(\myexu/_1323_ ), .ZN(\myexu/_0231_ ) );
INV_X1 \myexu/_4337_ ( .A(\myexu/_0387_ ), .ZN(\myexu/_1324_ ) );
NOR2_X1 \myexu/_4338_ ( .A1(\myexu/_0727_ ), .A2(\myexu/_2473_ ), .ZN(\myexu/_1325_ ) );
INV_X1 \myexu/_4339_ ( .A(\myexu/_1325_ ), .ZN(\myexu/_1326_ ) );
OAI21_X1 \myexu/_4340_ ( .A(\myexu/_1326_ ), .B1(\myexu/_1304_ ), .B2(\myexu/_1306_ ), .ZN(\myexu/_1327_ ) );
XNOR2_X1 \myexu/_4341_ ( .A(\myexu/_2442_ ), .B(\myexu/_2474_ ), .ZN(\myexu/_1328_ ) );
AOI21_X1 \myexu/_4342_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1327_ ), .B2(\myexu/_1328_ ), .ZN(\myexu/_1329_ ) );
OAI21_X1 \myexu/_4343_ ( .A(\myexu/_1329_ ), .B1(\myexu/_1327_ ), .B2(\myexu/_1328_ ), .ZN(\myexu/_1330_ ) );
NOR2_X1 \myexu/_4344_ ( .A1(\myexu/_0309_ ), .A2(\myexu/_2274_ ), .ZN(\myexu/_1331_ ) );
AND2_X1 \myexu/_4345_ ( .A1(\myexu/_0309_ ), .A2(\myexu/_2274_ ), .ZN(\myexu/_1332_ ) );
NOR3_X1 \myexu/_4346_ ( .A1(\myexu/_1312_ ), .A2(\myexu/_1331_ ), .A3(\myexu/_1332_ ), .ZN(\myexu/_1333_ ) );
NOR2_X1 \myexu/_4347_ ( .A1(\myexu/_1333_ ), .A2(\myexu/_1332_ ), .ZN(\myexu/_1334_ ) );
XOR2_X1 \myexu/_4348_ ( .A(\myexu/_0310_ ), .B(\myexu/_2275_ ), .Z(\myexu/_1335_ ) );
XNOR2_X1 \myexu/_4349_ ( .A(\myexu/_1334_ ), .B(\myexu/_1335_ ), .ZN(\myexu/_1336_ ) );
AOI22_X1 \myexu/_4350_ ( .A1(\myexu/_1336_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0310_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1337_ ) );
AOI21_X1 \myexu/_4351_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1330_ ), .B2(\myexu/_1337_ ), .ZN(\myexu/_1338_ ) );
AND2_X1 \myexu/_4352_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0049_ ), .ZN(\myexu/_1339_ ) );
NOR3_X1 \myexu/_4353_ ( .A1(\myexu/_1338_ ), .A2(\myexu/_1267_ ), .A3(\myexu/_1339_ ), .ZN(\myexu/_1340_ ) );
NAND3_X1 \myexu/_4354_ ( .A1(\myexu/_1319_ ), .A2(\myexu/_2274_ ), .A3(\myexu/_1320_ ), .ZN(\myexu/_1341_ ) );
XNOR2_X1 \myexu/_4355_ ( .A(\myexu/_1341_ ), .B(\myexu/_2275_ ), .ZN(\myexu/_1342_ ) );
OAI21_X1 \myexu/_4356_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1342_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_1343_ ) );
OAI21_X1 \myexu/_4357_ ( .A(\myexu/_1324_ ), .B1(\myexu/_1340_ ), .B2(\myexu/_1343_ ), .ZN(\myexu/_1344_ ) );
MUX2_X1 \myexu/_4358_ ( .A(\myexu/_2409_ ), .B(\myexu/_1344_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0232_ ) );
NAND3_X1 \myexu/_4359_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_1963_ ), .A3(\myexu/_2507_ ), .ZN(\myexu/_1345_ ) );
AND2_X1 \myexu/_4360_ ( .A1(\myexu/_1305_ ), .A2(\myexu/_1328_ ), .ZN(\myexu/_1346_ ) );
NAND2_X1 \myexu/_4361_ ( .A1(\myexu/_1303_ ), .A2(\myexu/_1346_ ), .ZN(\myexu/_1347_ ) );
NOR2_X1 \myexu/_4362_ ( .A1(\myexu/_1249_ ), .A2(\myexu/_1347_ ), .ZN(\myexu/_1348_ ) );
OAI21_X1 \myexu/_4363_ ( .A(\myexu/_1348_ ), .B1(\myexu/_1143_ ), .B2(\myexu/_1149_ ), .ZN(\myexu/_1349_ ) );
NAND2_X1 \myexu/_4364_ ( .A1(\myexu/_1328_ ), .A2(\myexu/_1325_ ), .ZN(\myexu/_1350_ ) );
OAI221_X1 \myexu/_4365_ ( .A(\myexu/_1350_ ), .B1(\myexu/_0384_ ), .B2(\myexu/_2474_ ), .C1(\myexu/_1248_ ), .C2(\myexu/_1347_ ), .ZN(\myexu/_1351_ ) );
AOI21_X1 \myexu/_4366_ ( .A(\myexu/_1351_ ), .B1(\myexu/_1302_ ), .B2(\myexu/_1346_ ), .ZN(\myexu/_1352_ ) );
NAND2_X2 \myexu/_4367_ ( .A1(\myexu/_1349_ ), .A2(\myexu/_1352_ ), .ZN(\myexu/_1353_ ) );
XNOR2_X1 \myexu/_4368_ ( .A(\myexu/_2443_ ), .B(\myexu/_2475_ ), .ZN(\myexu/_1354_ ) );
AND2_X1 \myexu/_4369_ ( .A1(\myexu/_1353_ ), .A2(\myexu/_1354_ ), .ZN(\myexu/_1355_ ) );
OAI21_X1 \myexu/_4370_ ( .A(\myexu/_0834_ ), .B1(\myexu/_1353_ ), .B2(\myexu/_1354_ ), .ZN(\myexu/_1356_ ) );
OR2_X1 \myexu/_4371_ ( .A1(\myexu/_1355_ ), .A2(\myexu/_1356_ ), .ZN(\myexu/_1357_ ) );
AND2_X1 \myexu/_4372_ ( .A1(\myexu/_1313_ ), .A2(\myexu/_1335_ ), .ZN(\myexu/_1358_ ) );
NAND3_X1 \myexu/_4373_ ( .A1(\myexu/_1358_ ), .A2(\myexu/_1261_ ), .A3(\myexu/_1289_ ), .ZN(\myexu/_1359_ ) );
AOI21_X2 \myexu/_4374_ ( .A(\myexu/_1359_ ), .B1(\myexu/_1255_ ), .B2(\myexu/_1259_ ), .ZN(\myexu/_1360_ ) );
AND4_X1 \myexu/_4375_ ( .A1(\myexu/_1310_ ), .A2(\myexu/_1313_ ), .A3(\myexu/_1335_ ), .A4(\myexu/_1311_ ), .ZN(\myexu/_1361_ ) );
AND2_X1 \myexu/_4376_ ( .A1(\myexu/_0310_ ), .A2(\myexu/_2275_ ), .ZN(\myexu/_1362_ ) );
AND2_X1 \myexu/_4377_ ( .A1(\myexu/_1335_ ), .A2(\myexu/_1332_ ), .ZN(\myexu/_1363_ ) );
OR3_X1 \myexu/_4378_ ( .A1(\myexu/_1361_ ), .A2(\myexu/_1362_ ), .A3(\myexu/_1363_ ), .ZN(\myexu/_1364_ ) );
OR2_X1 \myexu/_4379_ ( .A1(\myexu/_1360_ ), .A2(\myexu/_1364_ ), .ZN(\myexu/_1365_ ) );
XOR2_X1 \myexu/_4380_ ( .A(\myexu/_0311_ ), .B(\myexu/_2276_ ), .Z(\myexu/_1366_ ) );
XOR2_X1 \myexu/_4381_ ( .A(\myexu/_1365_ ), .B(\myexu/_1366_ ), .Z(\myexu/_1367_ ) );
AOI22_X1 \myexu/_4382_ ( .A1(\myexu/_1367_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0311_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1368_ ) );
AOI21_X1 \myexu/_4383_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1357_ ), .B2(\myexu/_1368_ ), .ZN(\myexu/_1369_ ) );
AND2_X1 \myexu/_4384_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0050_ ), .ZN(\myexu/_1370_ ) );
NOR3_X1 \myexu/_4385_ ( .A1(\myexu/_1369_ ), .A2(\myexu/_1267_ ), .A3(\myexu/_1370_ ), .ZN(\myexu/_1371_ ) );
AND2_X1 \myexu/_4386_ ( .A1(\myexu/_2274_ ), .A2(\myexu/_2275_ ), .ZN(\myexu/_1372_ ) );
NAND3_X1 \myexu/_4387_ ( .A1(\myexu/_1319_ ), .A2(\myexu/_1320_ ), .A3(\myexu/_1372_ ), .ZN(\myexu/_1373_ ) );
XNOR2_X1 \myexu/_4388_ ( .A(\myexu/_1373_ ), .B(\myexu/_2276_ ), .ZN(\myexu/_1374_ ) );
OAI21_X1 \myexu/_4389_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1374_ ), .B2(\myexu/_0865_ ), .ZN(\myexu/_1375_ ) );
OAI21_X1 \myexu/_4390_ ( .A(\myexu/_1345_ ), .B1(\myexu/_1371_ ), .B2(\myexu/_1375_ ), .ZN(\myexu/_1376_ ) );
MUX2_X1 \myexu/_4391_ ( .A(\myexu/_2410_ ), .B(\myexu/_1376_ ), .S(\myexu/_0981_ ), .Z(\myexu/_0233_ ) );
OAI21_X1 \myexu/_4392_ ( .A(\myexu/_2411_ ), .B1(\myexu/_1999_ ), .B2(fanout_net_5 ), .ZN(\myexu/_1377_ ) );
XNOR2_X1 \myexu/_4393_ ( .A(\myexu/_2444_ ), .B(\myexu/_2476_ ), .ZN(\myexu/_1378_ ) );
AND2_X1 \myexu/_4394_ ( .A1(\myexu/_1354_ ), .A2(\myexu/_1378_ ), .ZN(\myexu/_1379_ ) );
AND2_X1 \myexu/_4395_ ( .A1(\myexu/_1353_ ), .A2(\myexu/_1379_ ), .ZN(\myexu/_1380_ ) );
NOR2_X1 \myexu/_4396_ ( .A1(\myexu/_0392_ ), .A2(\myexu/_2475_ ), .ZN(\myexu/_1381_ ) );
AND2_X1 \myexu/_4397_ ( .A1(\myexu/_1378_ ), .A2(\myexu/_1381_ ), .ZN(\myexu/_1382_ ) );
INV_X1 \myexu/_4398_ ( .A(\myexu/_1382_ ), .ZN(\myexu/_1383_ ) );
NAND2_X1 \myexu/_4399_ ( .A1(\myexu/_1383_ ), .A2(\myexu/_0834_ ), .ZN(\myexu/_1384_ ) );
OR2_X1 \myexu/_4400_ ( .A1(\myexu/_1380_ ), .A2(\myexu/_1384_ ), .ZN(\myexu/_1385_ ) );
NOR3_X1 \myexu/_4401_ ( .A1(\myexu/_1355_ ), .A2(\myexu/_1381_ ), .A3(\myexu/_1378_ ), .ZN(\myexu/_1386_ ) );
OR2_X1 \myexu/_4402_ ( .A1(\myexu/_1385_ ), .A2(\myexu/_1386_ ), .ZN(\myexu/_1387_ ) );
OAI21_X1 \myexu/_4403_ ( .A(\myexu/_1366_ ), .B1(\myexu/_1360_ ), .B2(\myexu/_1364_ ), .ZN(\myexu/_1388_ ) );
NAND2_X1 \myexu/_4404_ ( .A1(\myexu/_0311_ ), .A2(\myexu/_2276_ ), .ZN(\myexu/_1389_ ) );
AND2_X1 \myexu/_4405_ ( .A1(\myexu/_1388_ ), .A2(\myexu/_1389_ ), .ZN(\myexu/_1390_ ) );
AND2_X1 \myexu/_4406_ ( .A1(\myexu/_0312_ ), .A2(\myexu/_2277_ ), .ZN(\myexu/_1391_ ) );
NOR2_X1 \myexu/_4407_ ( .A1(\myexu/_0312_ ), .A2(\myexu/_2277_ ), .ZN(\myexu/_1392_ ) );
NOR2_X1 \myexu/_4408_ ( .A1(\myexu/_1391_ ), .A2(\myexu/_1392_ ), .ZN(\myexu/_1393_ ) );
XNOR2_X1 \myexu/_4409_ ( .A(\myexu/_1390_ ), .B(\myexu/_1393_ ), .ZN(\myexu/_1394_ ) );
AOI22_X1 \myexu/_4410_ ( .A1(\myexu/_1394_ ), .A2(\myexu/_0853_ ), .B1(\myexu/_0312_ ), .B2(\myexu/_0854_ ), .ZN(\myexu/_1395_ ) );
AOI21_X1 \myexu/_4411_ ( .A(\myexu/_0845_ ), .B1(\myexu/_1387_ ), .B2(\myexu/_1395_ ), .ZN(\myexu/_1396_ ) );
AND2_X1 \myexu/_4412_ ( .A1(\myexu/_0792_ ), .A2(\myexu/_0051_ ), .ZN(\myexu/_1397_ ) );
NOR3_X1 \myexu/_4413_ ( .A1(\myexu/_1396_ ), .A2(\myexu/_0862_ ), .A3(\myexu/_1397_ ), .ZN(\myexu/_1398_ ) );
INV_X1 \myexu/_4414_ ( .A(\myexu/_2276_ ), .ZN(\myexu/_1399_ ) );
NOR2_X1 \myexu/_4415_ ( .A1(\myexu/_1373_ ), .A2(\myexu/_1399_ ), .ZN(\myexu/_1400_ ) );
XNOR2_X1 \myexu/_4416_ ( .A(\myexu/_1400_ ), .B(\myexu/_0406_ ), .ZN(\myexu/_1401_ ) );
OAI21_X1 \myexu/_4417_ ( .A(\myexu/_0931_ ), .B1(\myexu/_1401_ ), .B2(\myexu/_0866_ ), .ZN(\myexu/_1402_ ) );
OAI221_X1 \myexu/_4418_ ( .A(\myexu/_1377_ ), .B1(\myexu/_0401_ ), .B2(\myexu/_0844_ ), .C1(\myexu/_1398_ ), .C2(\myexu/_1402_ ), .ZN(\myexu/_0234_ ) );
NAND3_X1 \myexu/_4419_ ( .A1(\myexu/_2058_ ), .A2(\myexu/_1963_ ), .A3(\myexu/_2509_ ), .ZN(\myexu/_1403_ ) );
AOI21_X1 \myexu/_4420_ ( .A(\myexu/_1382_ ), .B1(\myexu/_2444_ ), .B2(\myexu/_0405_ ), .ZN(\myexu/_1404_ ) );
INV_X1 \myexu/_4421_ ( .A(\myexu/_1404_ ), .ZN(\myexu/_1405_ ) );
AOI21_X4 \myexu/_4422_ ( .A(\myexu/_1405_ ), .B1(\myexu/_1353_ ), .B2(\myexu/_1379_ ), .ZN(\myexu/_1406_ ) );
XNOR2_X1 \myexu/_4423_ ( .A(\myexu/_2445_ ), .B(\myexu/_2477_ ), .ZN(\myexu/_1407_ ) );
INV_X1 \myexu/_4424_ ( .A(\myexu/_1407_ ), .ZN(\myexu/_1408_ ) );
AOI21_X1 \myexu/_4425_ ( .A(\myexu/_0913_ ), .B1(\myexu/_1406_ ), .B2(\myexu/_1408_ ), .ZN(\myexu/_1409_ ) );
OAI21_X1 \myexu/_4426_ ( .A(\myexu/_1409_ ), .B1(\myexu/_1406_ ), .B2(\myexu/_1408_ ), .ZN(\myexu/_1410_ ) );
NOR3_X1 \myexu/_4427_ ( .A1(\myexu/_1391_ ), .A2(\myexu/_1392_ ), .A3(\myexu/_1389_ ), .ZN(\myexu/_1411_ ) );
OR2_X1 \myexu/_4428_ ( .A1(\myexu/_1411_ ), .A2(\myexu/_1391_ ), .ZN(\myexu/_1412_ ) );
AND2_X1 \myexu/_4429_ ( .A1(\myexu/_1366_ ), .A2(\myexu/_1393_ ), .ZN(\myexu/_1413_ ) );
AOI21_X1 \myexu/_4430_ ( .A(\myexu/_1412_ ), .B1(\myexu/_1365_ ), .B2(\myexu/_1413_ ), .ZN(\myexu/_1414_ ) );
XOR2_X1 \myexu/_4431_ ( .A(\myexu/_0313_ ), .B(\myexu/_2278_ ), .Z(\myexu/_1415_ ) );
XNOR2_X1 \myexu/_4432_ ( .A(\myexu/_1414_ ), .B(\myexu/_1415_ ), .ZN(\myexu/_1416_ ) );
AOI22_X1 \myexu/_4433_ ( .A1(\myexu/_1416_ ), .A2(\myexu/_0827_ ), .B1(\myexu/_0313_ ), .B2(\myexu/_0828_ ), .ZN(\myexu/_1417_ ) );
AOI21_X1 \myexu/_4434_ ( .A(\myexu/_0640_ ), .B1(\myexu/_1410_ ), .B2(\myexu/_1417_ ), .ZN(\myexu/_1418_ ) );
AND2_X1 \myexu/_4435_ ( .A1(\myexu/_0885_ ), .A2(\myexu/_0052_ ), .ZN(\myexu/_1419_ ) );
NOR3_X1 \myexu/_4436_ ( .A1(\myexu/_1418_ ), .A2(\myexu/_1267_ ), .A3(\myexu/_1419_ ), .ZN(\myexu/_1420_ ) );
AND4_X1 \myexu/_4437_ ( .A1(\myexu/_2276_ ), .A2(\myexu/_1320_ ), .A3(\myexu/_2277_ ), .A4(\myexu/_1372_ ), .ZN(\myexu/_1421_ ) );
AND2_X1 \myexu/_4438_ ( .A1(\myexu/_1319_ ), .A2(\myexu/_1421_ ), .ZN(\myexu/_1422_ ) );
INV_X1 \myexu/_4439_ ( .A(\myexu/_2278_ ), .ZN(\myexu/_1423_ ) );
XNOR2_X1 \myexu/_4440_ ( .A(\myexu/_1422_ ), .B(\myexu/_1423_ ), .ZN(\myexu/_1424_ ) );
OAI21_X1 \myexu/_4441_ ( .A(\myexu/_0819_ ), .B1(\myexu/_1424_ ), .B2(\myexu/_0796_ ), .ZN(\myexu/_1425_ ) );
OAI21_X1 \myexu/_4442_ ( .A(\myexu/_1403_ ), .B1(\myexu/_1420_ ), .B2(\myexu/_1425_ ), .ZN(\myexu/_1426_ ) );
MUX2_X1 \myexu/_4443_ ( .A(\myexu/_2412_ ), .B(\myexu/_1426_ ), .S(\myexu/_2012_ ), .Z(\myexu/_0235_ ) );
NOR2_X4 \myexu/_4444_ ( .A1(\myexu/_1406_ ), .A2(\myexu/_1408_ ), .ZN(\myexu/_1427_ ) );
NOR2_X1 \myexu/_4445_ ( .A1(\myexu/_0410_ ), .A2(\myexu/_2477_ ), .ZN(\myexu/_1428_ ) );
OR2_X1 \myexu/_4446_ ( .A1(\myexu/_1427_ ), .A2(\myexu/_1428_ ), .ZN(\myexu/_1429_ ) );
XNOR2_X1 \myexu/_4447_ ( .A(\myexu/_2446_ ), .B(\myexu/_2478_ ), .ZN(\myexu/_1430_ ) );
AOI21_X1 \myexu/_4448_ ( .A(\myexu/_0773_ ), .B1(\myexu/_1429_ ), .B2(\myexu/_1430_ ), .ZN(\myexu/_1431_ ) );
OAI21_X1 \myexu/_4449_ ( .A(\myexu/_1431_ ), .B1(\myexu/_1429_ ), .B2(\myexu/_1430_ ), .ZN(\myexu/_1432_ ) );
NOR2_X1 \myexu/_4450_ ( .A1(\myexu/_0313_ ), .A2(\myexu/_2278_ ), .ZN(\myexu/_1433_ ) );
AND2_X1 \myexu/_4451_ ( .A1(\myexu/_0313_ ), .A2(\myexu/_2278_ ), .ZN(\myexu/_1434_ ) );
NOR3_X1 \myexu/_4452_ ( .A1(\myexu/_1414_ ), .A2(\myexu/_1433_ ), .A3(\myexu/_1434_ ), .ZN(\myexu/_1435_ ) );
NOR2_X1 \myexu/_4453_ ( .A1(\myexu/_1435_ ), .A2(\myexu/_1434_ ), .ZN(\myexu/_1436_ ) );
XOR2_X1 \myexu/_4454_ ( .A(\myexu/_0314_ ), .B(\myexu/_2279_ ), .Z(\myexu/_1437_ ) );
XNOR2_X1 \myexu/_4455_ ( .A(\myexu/_1436_ ), .B(\myexu/_1437_ ), .ZN(\myexu/_1438_ ) );
AOI22_X1 \myexu/_4456_ ( .A1(\myexu/_1438_ ), .A2(\myexu/_0780_ ), .B1(\myexu/_0314_ ), .B2(\myexu/_0778_ ), .ZN(\myexu/_1439_ ) );
AOI21_X1 \myexu/_4457_ ( .A(\myexu/_0639_ ), .B1(\myexu/_1432_ ), .B2(\myexu/_1439_ ), .ZN(\myexu/_1440_ ) );
AND2_X1 \myexu/_4458_ ( .A1(\myexu/_0791_ ), .A2(\myexu/_0053_ ), .ZN(\myexu/_1441_ ) );
OR3_X1 \myexu/_4459_ ( .A1(\myexu/_1440_ ), .A2(\myexu/_0786_ ), .A3(\myexu/_1441_ ), .ZN(\myexu/_1442_ ) );
NAND3_X1 \myexu/_4460_ ( .A1(\myexu/_1319_ ), .A2(\myexu/_2278_ ), .A3(\myexu/_1421_ ), .ZN(\myexu/_1443_ ) );
XNOR2_X1 \myexu/_4461_ ( .A(\myexu/_1443_ ), .B(\myexu/_2279_ ), .ZN(\myexu/_1444_ ) );
OR2_X1 \myexu/_4462_ ( .A1(\myexu/_1444_ ), .A2(\myexu/_0796_ ), .ZN(\myexu/_1445_ ) );
NAND3_X1 \myexu/_4463_ ( .A1(\myexu/_1442_ ), .A2(\myexu/_2140_ ), .A3(\myexu/_1445_ ), .ZN(\myexu/_1446_ ) );
INV_X1 \myexu/_4464_ ( .A(\myexu/_2510_ ), .ZN(\myexu/_1447_ ) );
OAI21_X1 \myexu/_4465_ ( .A(\myexu/_1446_ ), .B1(\myexu/_1447_ ), .B2(\myexu/_2140_ ), .ZN(\myexu/_1448_ ) );
MUX2_X1 \myexu/_4466_ ( .A(\myexu/_2413_ ), .B(\myexu/_1448_ ), .S(\myexu/_2012_ ), .Z(\myexu/_0236_ ) );
NOR2_X1 \myexu/_4467_ ( .A1(\myexu/_0418_ ), .A2(\myexu/_2446_ ), .ZN(\myexu/_1449_ ) );
INV_X2 \myexu/_4468_ ( .A(\myexu/_1427_ ), .ZN(\myexu/_1450_ ) );
AOI21_X1 \myexu/_4469_ ( .A(\myexu/_1428_ ), .B1(\myexu/_2446_ ), .B2(\myexu/_0418_ ), .ZN(\myexu/_1451_ ) );
AOI21_X4 \myexu/_4470_ ( .A(\myexu/_1449_ ), .B1(\myexu/_1450_ ), .B2(\myexu/_1451_ ), .ZN(\myexu/_1452_ ) );
XNOR2_X1 \myexu/_4471_ ( .A(\myexu/_2447_ ), .B(\myexu/_2479_ ), .ZN(\myexu/_1453_ ) );
AND2_X1 \myexu/_4472_ ( .A1(\myexu/_1452_ ), .A2(\myexu/_1453_ ), .ZN(\myexu/_1454_ ) );
OAI21_X1 \myexu/_4473_ ( .A(\myexu/_0834_ ), .B1(\myexu/_1452_ ), .B2(\myexu/_1453_ ), .ZN(\myexu/_1455_ ) );
NOR2_X1 \myexu/_4474_ ( .A1(\myexu/_1454_ ), .A2(\myexu/_1455_ ), .ZN(\myexu/_1456_ ) );
AND2_X1 \myexu/_4475_ ( .A1(\myexu/_1415_ ), .A2(\myexu/_1437_ ), .ZN(\myexu/_1457_ ) );
OAI211_X2 \myexu/_4476_ ( .A(\myexu/_1413_ ), .B(\myexu/_1457_ ), .C1(\myexu/_1360_ ), .C2(\myexu/_1364_ ), .ZN(\myexu/_1458_ ) );
AND2_X1 \myexu/_4477_ ( .A1(\myexu/_1437_ ), .A2(\myexu/_1434_ ), .ZN(\myexu/_1459_ ) );
AOI221_X4 \myexu/_4478_ ( .A(\myexu/_1459_ ), .B1(\myexu/_0314_ ), .B2(\myexu/_2279_ ), .C1(\myexu/_1412_ ), .C2(\myexu/_1457_ ), .ZN(\myexu/_1460_ ) );
NAND2_X1 \myexu/_4479_ ( .A1(\myexu/_1458_ ), .A2(\myexu/_1460_ ), .ZN(\myexu/_1461_ ) );
XOR2_X1 \myexu/_4480_ ( .A(\myexu/_0315_ ), .B(\myexu/_2280_ ), .Z(\myexu/_1462_ ) );
INV_X1 \myexu/_4481_ ( .A(\myexu/_1462_ ), .ZN(\myexu/_1463_ ) );
XNOR2_X1 \myexu/_4482_ ( .A(\myexu/_1461_ ), .B(\myexu/_1463_ ), .ZN(\myexu/_1464_ ) );
INV_X1 \myexu/_4483_ ( .A(\myexu/_1464_ ), .ZN(\myexu/_1465_ ) );
OAI22_X1 \myexu/_4484_ ( .A1(\myexu/_1465_ ), .A2(\myexu/_0805_ ), .B1(\myexu/_0431_ ), .B2(\myexu/_0806_ ), .ZN(\myexu/_1466_ ) );
OAI21_X1 \myexu/_4485_ ( .A(\myexu/_0800_ ), .B1(\myexu/_1456_ ), .B2(\myexu/_1466_ ), .ZN(\myexu/_1467_ ) );
OAI21_X1 \myexu/_4486_ ( .A(\myexu/_0054_ ), .B1(\myexu/_0789_ ), .B2(\myexu/_0639_ ), .ZN(\myexu/_1468_ ) );
NAND3_X1 \myexu/_4487_ ( .A1(\myexu/_1467_ ), .A2(\myexu/_0795_ ), .A3(\myexu/_1468_ ), .ZN(\myexu/_1469_ ) );
AND3_X1 \myexu/_4488_ ( .A1(\myexu/_1422_ ), .A2(\myexu/_2278_ ), .A3(\myexu/_2279_ ), .ZN(\myexu/_1470_ ) );
XNOR2_X1 \myexu/_4489_ ( .A(\myexu/_1470_ ), .B(\myexu/_2280_ ), .ZN(\myexu/_1471_ ) );
NAND2_X1 \myexu/_4490_ ( .A1(\myexu/_1471_ ), .A2(\myexu/_0786_ ), .ZN(\myexu/_1472_ ) );
AND3_X1 \myexu/_4491_ ( .A1(\myexu/_1469_ ), .A2(\myexu/_2131_ ), .A3(\myexu/_1472_ ), .ZN(\myexu/_1473_ ) );
OR2_X1 \myexu/_4492_ ( .A1(\myexu/_1473_ ), .A2(\myexu/_0436_ ), .ZN(\myexu/_1474_ ) );
MUX2_X1 \myexu/_4493_ ( .A(\myexu/_2414_ ), .B(\myexu/_1474_ ), .S(\myexu/_2012_ ), .Z(\myexu/_0237_ ) );
NOR2_X1 \myexu/_4494_ ( .A1(\myexu/_0642_ ), .A2(\myexu/_2479_ ), .ZN(\myexu/_1475_ ) );
XNOR2_X1 \myexu/_4495_ ( .A(\myexu/_2448_ ), .B(\myexu/_2480_ ), .ZN(\myexu/_1476_ ) );
OR3_X4 \myexu/_4496_ ( .A1(\myexu/_1454_ ), .A2(\myexu/_1475_ ), .A3(\myexu/_1476_ ), .ZN(\myexu/_1477_ ) );
AND2_X1 \myexu/_4497_ ( .A1(\myexu/_1476_ ), .A2(\myexu/_1475_ ), .ZN(\myexu/_1478_ ) );
AND2_X1 \myexu/_4498_ ( .A1(\myexu/_1453_ ), .A2(\myexu/_1476_ ), .ZN(\myexu/_1479_ ) );
AOI211_X4 \myexu/_4499_ ( .A(\myexu/_0772_ ), .B(\myexu/_1478_ ), .C1(\myexu/_1452_ ), .C2(\myexu/_1479_ ), .ZN(\myexu/_1480_ ) );
AND2_X1 \myexu/_4500_ ( .A1(\myexu/_1477_ ), .A2(\myexu/_1480_ ), .ZN(\myexu/_1481_ ) );
NAND2_X1 \myexu/_4501_ ( .A1(\myexu/_1461_ ), .A2(\myexu/_1462_ ), .ZN(\myexu/_1482_ ) );
NAND2_X1 \myexu/_4502_ ( .A1(\myexu/_0315_ ), .A2(\myexu/_2280_ ), .ZN(\myexu/_1483_ ) );
NAND2_X1 \myexu/_4503_ ( .A1(\myexu/_1482_ ), .A2(\myexu/_1483_ ), .ZN(\myexu/_1484_ ) );
XNOR2_X1 \myexu/_4504_ ( .A(\myexu/_0316_ ), .B(\myexu/_2281_ ), .ZN(\myexu/_1485_ ) );
XNOR2_X1 \myexu/_4505_ ( .A(\myexu/_1484_ ), .B(\myexu/_1485_ ), .ZN(\myexu/_1486_ ) );
AND2_X1 \myexu/_4506_ ( .A1(\myexu/_1486_ ), .A2(\myexu/_0780_ ), .ZN(\myexu/_1487_ ) );
AND3_X1 \myexu/_4507_ ( .A1(\myexu/_0776_ ), .A2(\myexu/_0777_ ), .A3(\myexu/_0316_ ), .ZN(\myexu/_1488_ ) );
OR2_X1 \myexu/_4508_ ( .A1(\myexu/_1487_ ), .A2(\myexu/_1488_ ), .ZN(\myexu/_1489_ ) );
OAI21_X1 \myexu/_4509_ ( .A(\myexu/_0800_ ), .B1(\myexu/_1481_ ), .B2(\myexu/_1489_ ), .ZN(\myexu/_1490_ ) );
AOI21_X1 \myexu/_4510_ ( .A(\myexu/_0785_ ), .B1(\myexu/_0791_ ), .B2(\myexu/_0055_ ), .ZN(\myexu/_1491_ ) );
NAND2_X1 \myexu/_4511_ ( .A1(\myexu/_1470_ ), .A2(\myexu/_2280_ ), .ZN(\myexu/_1492_ ) );
XNOR2_X1 \myexu/_4512_ ( .A(\myexu/_1492_ ), .B(\myexu/_0441_ ), .ZN(\myexu/_1493_ ) );
AOI22_X1 \myexu/_4513_ ( .A1(\myexu/_1490_ ), .A2(\myexu/_1491_ ), .B1(\myexu/_0786_ ), .B2(\myexu/_1493_ ), .ZN(\myexu/_1494_ ) );
MUX2_X1 \myexu/_4514_ ( .A(\myexu/_2512_ ), .B(\myexu/_1494_ ), .S(\myexu/_2131_ ), .Z(\myexu/_1495_ ) );
MUX2_X1 \myexu/_4515_ ( .A(\myexu/_2415_ ), .B(\myexu/_1495_ ), .S(\myexu/_2012_ ), .Z(\myexu/_0238_ ) );
AND3_X4 \myexu/_4516_ ( .A1(\myexu/_1117_ ), .A2(\myexu/_2265_ ), .A3(\myexu/_2266_ ), .ZN(\myexu/_1496_ ) );
AND3_X1 \myexu/_4517_ ( .A1(\myexu/_1496_ ), .A2(\myexu/_2267_ ), .A3(\myexu/_2268_ ), .ZN(\myexu/_1497_ ) );
AND2_X1 \myexu/_4518_ ( .A1(\myexu/_1497_ ), .A2(\myexu/_2269_ ), .ZN(\myexu/_1498_ ) );
AND3_X1 \myexu/_4519_ ( .A1(\myexu/_1498_ ), .A2(\myexu/_2270_ ), .A3(\myexu/_2272_ ), .ZN(\myexu/_1499_ ) );
AND2_X1 \myexu/_4520_ ( .A1(\myexu/_1499_ ), .A2(\myexu/_2273_ ), .ZN(\myexu/_1500_ ) );
AND2_X1 \myexu/_4521_ ( .A1(\myexu/_1500_ ), .A2(\myexu/_2274_ ), .ZN(\myexu/_1501_ ) );
AND3_X1 \myexu/_4522_ ( .A1(\myexu/_1501_ ), .A2(\myexu/_2275_ ), .A3(\myexu/_2276_ ), .ZN(\myexu/_1502_ ) );
AND3_X1 \myexu/_4523_ ( .A1(\myexu/_1502_ ), .A2(\myexu/_2277_ ), .A3(\myexu/_2278_ ), .ZN(\myexu/_1503_ ) );
AND3_X2 \myexu/_4524_ ( .A1(\myexu/_1503_ ), .A2(\myexu/_2279_ ), .A3(\myexu/_2280_ ), .ZN(\myexu/_1504_ ) );
AND2_X1 \myexu/_4525_ ( .A1(\myexu/_1504_ ), .A2(\myexu/_2281_ ), .ZN(\myexu/_1505_ ) );
XOR2_X1 \myexu/_4526_ ( .A(\myexu/_1505_ ), .B(\myexu/_2283_ ), .Z(\myexu/_1506_ ) );
NOR2_X1 \myexu/_4527_ ( .A1(\myexu/_1506_ ), .A2(\myexu/_0795_ ), .ZN(\myexu/_1507_ ) );
AOI21_X1 \myexu/_4528_ ( .A(\myexu/_1478_ ), .B1(\myexu/_2448_ ), .B2(\myexu/_0439_ ), .ZN(\myexu/_1508_ ) );
INV_X1 \myexu/_4529_ ( .A(\myexu/_1508_ ), .ZN(\myexu/_1509_ ) );
AOI21_X4 \myexu/_4530_ ( .A(\myexu/_1509_ ), .B1(\myexu/_1452_ ), .B2(\myexu/_1479_ ), .ZN(\myexu/_1510_ ) );
XNOR2_X1 \myexu/_4531_ ( .A(\myexu/_2450_ ), .B(\myexu/_2482_ ), .ZN(\myexu/_1511_ ) );
INV_X1 \myexu/_4532_ ( .A(\myexu/_1511_ ), .ZN(\myexu/_1512_ ) );
NOR2_X2 \myexu/_4533_ ( .A1(\myexu/_1510_ ), .A2(\myexu/_1512_ ), .ZN(\myexu/_1513_ ) );
INV_X1 \myexu/_4534_ ( .A(\myexu/_1513_ ), .ZN(\myexu/_1514_ ) );
AOI21_X1 \myexu/_4535_ ( .A(\myexu/_0773_ ), .B1(\myexu/_1510_ ), .B2(\myexu/_1512_ ), .ZN(\myexu/_1515_ ) );
AND2_X1 \myexu/_4536_ ( .A1(\myexu/_1514_ ), .A2(\myexu/_1515_ ), .ZN(\myexu/_1516_ ) );
AOI211_X2 \myexu/_4537_ ( .A(\myexu/_1463_ ), .B(\myexu/_1485_ ), .C1(\myexu/_1458_ ), .C2(\myexu/_1460_ ), .ZN(\myexu/_1517_ ) );
AND2_X1 \myexu/_4538_ ( .A1(\myexu/_0316_ ), .A2(\myexu/_2281_ ), .ZN(\myexu/_1518_ ) );
NOR2_X1 \myexu/_4539_ ( .A1(\myexu/_1485_ ), .A2(\myexu/_1483_ ), .ZN(\myexu/_1519_ ) );
NOR3_X1 \myexu/_4540_ ( .A1(\myexu/_1517_ ), .A2(\myexu/_1518_ ), .A3(\myexu/_1519_ ), .ZN(\myexu/_1520_ ) );
XNOR2_X1 \myexu/_4541_ ( .A(\myexu/_0318_ ), .B(\myexu/_2283_ ), .ZN(\myexu/_1521_ ) );
XOR2_X1 \myexu/_4542_ ( .A(\myexu/_1520_ ), .B(\myexu/_1521_ ), .Z(\myexu/_1522_ ) );
NAND2_X1 \myexu/_4543_ ( .A1(\myexu/_1522_ ), .A2(\myexu/_0780_ ), .ZN(\myexu/_1523_ ) );
OAI21_X1 \myexu/_4544_ ( .A(\myexu/_1523_ ), .B1(\myexu/_0456_ ), .B2(\myexu/_0806_ ), .ZN(\myexu/_1524_ ) );
OAI21_X1 \myexu/_4545_ ( .A(\myexu/_0800_ ), .B1(\myexu/_1516_ ), .B2(\myexu/_1524_ ), .ZN(\myexu/_1525_ ) );
AOI21_X1 \myexu/_4546_ ( .A(\myexu/_0786_ ), .B1(\myexu/_0791_ ), .B2(\myexu/_0057_ ), .ZN(\myexu/_1526_ ) );
AOI21_X1 \myexu/_4547_ ( .A(\myexu/_1507_ ), .B1(\myexu/_1525_ ), .B2(\myexu/_1526_ ), .ZN(\myexu/_1527_ ) );
MUX2_X1 \myexu/_4548_ ( .A(\myexu/_2514_ ), .B(\myexu/_1527_ ), .S(\myexu/_2131_ ), .Z(\myexu/_1528_ ) );
MUX2_X1 \myexu/_4549_ ( .A(\myexu/_2417_ ), .B(\myexu/_1528_ ), .S(\myexu/_2012_ ), .Z(\myexu/_0239_ ) );
NOR2_X1 \myexu/_4550_ ( .A1(\myexu/_0755_ ), .A2(\myexu/_2482_ ), .ZN(\myexu/_1529_ ) );
XNOR2_X1 \myexu/_4551_ ( .A(\myexu/_2483_ ), .B(\myexu/_2451_ ), .ZN(\myexu/_1530_ ) );
OR3_X4 \myexu/_4552_ ( .A1(\myexu/_1513_ ), .A2(\myexu/_1529_ ), .A3(\myexu/_1530_ ), .ZN(\myexu/_1531_ ) );
OAI21_X1 \myexu/_4553_ ( .A(\myexu/_1530_ ), .B1(\myexu/_1513_ ), .B2(\myexu/_1529_ ), .ZN(\myexu/_1532_ ) );
NAND3_X1 \myexu/_4554_ ( .A1(\myexu/_1531_ ), .A2(\myexu/_0834_ ), .A3(\myexu/_1532_ ), .ZN(\myexu/_1533_ ) );
NOR2_X1 \myexu/_4555_ ( .A1(\myexu/_1520_ ), .A2(\myexu/_1521_ ), .ZN(\myexu/_1534_ ) );
AND2_X1 \myexu/_4556_ ( .A1(\myexu/_0318_ ), .A2(\myexu/_2283_ ), .ZN(\myexu/_1535_ ) );
NOR2_X1 \myexu/_4557_ ( .A1(\myexu/_1534_ ), .A2(\myexu/_1535_ ), .ZN(\myexu/_1536_ ) );
XNOR2_X1 \myexu/_4558_ ( .A(\myexu/_0319_ ), .B(\myexu/_2284_ ), .ZN(\myexu/_1537_ ) );
XOR2_X1 \myexu/_4559_ ( .A(\myexu/_1536_ ), .B(\myexu/_1537_ ), .Z(\myexu/_1538_ ) );
AOI22_X1 \myexu/_4560_ ( .A1(\myexu/_1538_ ), .A2(\myexu/_0780_ ), .B1(\myexu/_0319_ ), .B2(\myexu/_0778_ ), .ZN(\myexu/_1539_ ) );
AOI21_X1 \myexu/_4561_ ( .A(\myexu/_0639_ ), .B1(\myexu/_1533_ ), .B2(\myexu/_1539_ ), .ZN(\myexu/_1540_ ) );
AND2_X1 \myexu/_4562_ ( .A1(\myexu/_0791_ ), .A2(\myexu/_0058_ ), .ZN(\myexu/_1541_ ) );
NOR3_X1 \myexu/_4563_ ( .A1(\myexu/_1540_ ), .A2(\myexu/_0785_ ), .A3(\myexu/_1541_ ), .ZN(\myexu/_1542_ ) );
NAND3_X1 \myexu/_4564_ ( .A1(\myexu/_1504_ ), .A2(\myexu/_2281_ ), .A3(\myexu/_2283_ ), .ZN(\myexu/_1543_ ) );
INV_X1 \myexu/_4565_ ( .A(\myexu/_2284_ ), .ZN(\myexu/_1544_ ) );
XNOR2_X1 \myexu/_4566_ ( .A(\myexu/_1543_ ), .B(\myexu/_1544_ ), .ZN(\myexu/_1545_ ) );
AOI21_X1 \myexu/_4567_ ( .A(\myexu/_1542_ ), .B1(\myexu/_1267_ ), .B2(\myexu/_1545_ ), .ZN(\myexu/_1546_ ) );
MUX2_X2 \myexu/_4568_ ( .A(\myexu/_2515_ ), .B(\myexu/_1546_ ), .S(\myexu/_2131_ ), .Z(\myexu/_1547_ ) );
MUX2_X2 \myexu/_4569_ ( .A(\myexu/_2418_ ), .B(\myexu/_1547_ ), .S(\myexu/_2012_ ), .Z(\myexu/_0240_ ) );
NAND2_X1 \myexu/_4570_ ( .A1(\myexu/_1981_ ), .A2(\myexu/_2530_ ), .ZN(\myexu/_1548_ ) );
NOR2_X1 \myexu/_4571_ ( .A1(\myexu/_0816_ ), .A2(\myexu/_2528_ ), .ZN(\myexu/_1549_ ) );
NOR2_X2 \myexu/_4572_ ( .A1(\myexu/_1548_ ), .A2(\myexu/_1549_ ), .ZN(\myexu/_1550_ ) );
BUF_X8 \myexu/_4573_ ( .A(\myexu/_1550_ ), .Z(\myexu/_1551_ ) );
BUF_X8 \myexu/_4574_ ( .A(\myexu/_2030_ ), .Z(\myexu/_1552_ ) );
BUF_X4 \myexu/_4575_ ( .A(\myexu/_1267_ ), .Z(\myexu/_1553_ ) );
NAND3_X1 \myexu/_4576_ ( .A1(\myexu/_0761_ ), .A2(\myexu/_2118_ ), .A3(\myexu/_2108_ ), .ZN(\myexu/_1554_ ) );
AND2_X1 \myexu/_4577_ ( .A1(\myexu/_1407_ ), .A2(\myexu/_1430_ ), .ZN(\myexu/_1555_ ) );
AND2_X1 \myexu/_4578_ ( .A1(\myexu/_1379_ ), .A2(\myexu/_1555_ ), .ZN(\myexu/_1556_ ) );
AND3_X1 \myexu/_4579_ ( .A1(\myexu/_1479_ ), .A2(\myexu/_1511_ ), .A3(\myexu/_1530_ ), .ZN(\myexu/_1557_ ) );
AND3_X1 \myexu/_4580_ ( .A1(\myexu/_1348_ ), .A2(\myexu/_1556_ ), .A3(\myexu/_1557_ ), .ZN(\myexu/_1558_ ) );
OAI21_X1 \myexu/_4581_ ( .A(\myexu/_1558_ ), .B1(\myexu/_1143_ ), .B2(\myexu/_1149_ ), .ZN(\myexu/_1559_ ) );
AND2_X1 \myexu/_4582_ ( .A1(\myexu/_1557_ ), .A2(\myexu/_1556_ ), .ZN(\myexu/_1560_ ) );
INV_X1 \myexu/_4583_ ( .A(\myexu/_1560_ ), .ZN(\myexu/_1561_ ) );
OR2_X1 \myexu/_4584_ ( .A1(\myexu/_1352_ ), .A2(\myexu/_1561_ ), .ZN(\myexu/_1562_ ) );
NAND2_X1 \myexu/_4585_ ( .A1(\myexu/_1405_ ), .A2(\myexu/_1555_ ), .ZN(\myexu/_1563_ ) );
OAI21_X1 \myexu/_4586_ ( .A(\myexu/_1563_ ), .B1(\myexu/_1449_ ), .B2(\myexu/_1451_ ), .ZN(\myexu/_1564_ ) );
NAND2_X1 \myexu/_4587_ ( .A1(\myexu/_1564_ ), .A2(\myexu/_1557_ ), .ZN(\myexu/_1565_ ) );
NAND3_X1 \myexu/_4588_ ( .A1(\myexu/_1509_ ), .A2(\myexu/_1511_ ), .A3(\myexu/_1530_ ), .ZN(\myexu/_1566_ ) );
NOR2_X1 \myexu/_4589_ ( .A1(\myexu/_0465_ ), .A2(\myexu/_2483_ ), .ZN(\myexu/_1567_ ) );
AOI21_X1 \myexu/_4590_ ( .A(\myexu/_1567_ ), .B1(\myexu/_1530_ ), .B2(\myexu/_1529_ ), .ZN(\myexu/_1568_ ) );
AND4_X1 \myexu/_4591_ ( .A1(\myexu/_1562_ ), .A2(\myexu/_1565_ ), .A3(\myexu/_1566_ ), .A4(\myexu/_1568_ ), .ZN(\myexu/_1569_ ) );
AND2_X2 \myexu/_4592_ ( .A1(\myexu/_1559_ ), .A2(\myexu/_1569_ ), .ZN(\myexu/_1570_ ) );
NAND3_X1 \myexu/_4593_ ( .A1(\myexu/_1570_ ), .A2(\myexu/_2525_ ), .A3(\myexu/_0764_ ), .ZN(\myexu/_1571_ ) );
OR3_X2 \myexu/_4594_ ( .A1(\myexu/_1570_ ), .A2(\myexu/_2118_ ), .A3(\myexu/_0444_ ), .ZN(\myexu/_1572_ ) );
AND4_X1 \myexu/_4595_ ( .A1(\myexu/_0774_ ), .A2(\myexu/_0808_ ), .A3(\myexu/_0916_ ), .A4(\myexu/_0945_ ), .ZN(\myexu/_1573_ ) );
AND4_X1 \myexu/_4596_ ( .A1(\myexu/_0832_ ), .A2(\myexu/_0857_ ), .A3(\myexu/_0880_ ), .A4(\myexu/_0893_ ), .ZN(\myexu/_1574_ ) );
AND4_X1 \myexu/_4597_ ( .A1(\myexu/_1053_ ), .A2(\myexu/_1142_ ), .A3(\myexu/_1573_ ), .A4(\myexu/_1574_ ), .ZN(\myexu/_1575_ ) );
NAND3_X1 \myexu/_4598_ ( .A1(\myexu/_2107_ ), .A2(\myexu/_2112_ ), .A3(fanout_net_7 ), .ZN(\myexu/_1576_ ) );
NAND4_X1 \myexu/_4599_ ( .A1(\myexu/_1560_ ), .A2(\myexu/_1575_ ), .A3(\myexu/_1348_ ), .A4(\myexu/_1576_ ), .ZN(\myexu/_1577_ ) );
AND2_X1 \myexu/_4600_ ( .A1(\myexu/_1558_ ), .A2(\myexu/_1575_ ), .ZN(\myexu/_1578_ ) );
OAI21_X1 \myexu/_4601_ ( .A(\myexu/_1577_ ), .B1(\myexu/_1578_ ), .B2(\myexu/_0767_ ), .ZN(\myexu/_1579_ ) );
AND4_X2 \myexu/_4602_ ( .A1(\myexu/_1554_ ), .A2(\myexu/_1571_ ), .A3(\myexu/_1572_ ), .A4(\myexu/_1579_ ), .ZN(\myexu/_1580_ ) );
NOR3_X1 \myexu/_4603_ ( .A1(\myexu/_2113_ ), .A2(fanout_net_7 ), .A3(\myexu/_2524_ ), .ZN(\myexu/_1581_ ) );
NAND3_X1 \myexu/_4604_ ( .A1(\myexu/_0759_ ), .A2(\myexu/_0760_ ), .A3(\myexu/_1581_ ), .ZN(\myexu/_1582_ ) );
AND2_X4 \myexu/_4605_ ( .A1(\myexu/_1580_ ), .A2(\myexu/_1582_ ), .ZN(\myexu/_1583_ ) );
BUF_X16 \myexu/_4606_ ( .A(\myexu/_1583_ ), .Z(\myexu/_1584_ ) );
BUF_X4 \myexu/_4607_ ( .A(\myexu/_1584_ ), .Z(\myexu/_1585_ ) );
BUF_X2 \myexu/_4608_ ( .A(\myexu/_1585_ ), .Z(\myexu/_1586_ ) );
OR2_X1 \myexu/_4609_ ( .A1(\myexu/_1586_ ), .A2(\myexu/_2260_ ), .ZN(\myexu/_1587_ ) );
BUF_X4 \myexu/_4610_ ( .A(\myexu/_0762_ ), .Z(\myexu/_1588_ ) );
BUF_X4 \myexu/_4611_ ( .A(\myexu/_1588_ ), .Z(\myexu/_1589_ ) );
INV_X8 \myexu/_4612_ ( .A(\myexu/_1584_ ), .ZN(\myexu/_1590_ ) );
BUF_X4 \myexu/_4613_ ( .A(\myexu/_1590_ ), .Z(\myexu/_1591_ ) );
OAI211_X2 \myexu/_4614_ ( .A(\myexu/_1587_ ), .B(\myexu/_1589_ ), .C1(\myexu/_0781_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1592_ ) );
NAND2_X1 \myexu/_4615_ ( .A1(\myexu/_2491_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1593_ ) );
AOI21_X1 \myexu/_4616_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1592_ ), .B2(\myexu/_1593_ ), .ZN(\myexu/_1594_ ) );
NAND3_X1 \myexu/_4617_ ( .A1(\myexu/_0787_ ), .A2(\myexu/_2121_ ), .A3(\myexu/_0781_ ), .ZN(\myexu/_1595_ ) );
NAND2_X1 \myexu/_4618_ ( .A1(\myexu/_1595_ ), .A2(\myexu/_0440_ ), .ZN(\myexu/_1596_ ) );
OAI221_X1 \myexu/_4619_ ( .A(\myexu/_1551_ ), .B1(\myexu/_2491_ ), .B2(\myexu/_1552_ ), .C1(\myexu/_1594_ ), .C2(\myexu/_1596_ ), .ZN(\myexu/_1597_ ) );
BUF_X4 \myexu/_4620_ ( .A(\myexu/_1548_ ), .Z(\myexu/_1598_ ) );
BUF_X4 \myexu/_4621_ ( .A(\myexu/_1598_ ), .Z(\myexu/_1599_ ) );
BUF_X4 \myexu/_4622_ ( .A(\myexu/_1549_ ), .Z(\myexu/_1600_ ) );
BUF_X4 \myexu/_4623_ ( .A(\myexu/_1600_ ), .Z(\myexu/_1601_ ) );
OAI21_X1 \myexu/_4624_ ( .A(\myexu/_2292_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1602_ ) );
AOI21_X1 \myexu/_4625_ ( .A(fanout_net_5 ), .B1(\myexu/_1597_ ), .B2(\myexu/_1602_ ), .ZN(\myexu/_0110_ ) );
BUF_X4 \myexu/_4626_ ( .A(\myexu/_1550_ ), .Z(\myexu/_1603_ ) );
BUF_X4 \myexu/_4627_ ( .A(\myexu/_2030_ ), .Z(\myexu/_1604_ ) );
MUX2_X1 \myexu/_4628_ ( .A(\myexu/_2271_ ), .B(\myexu/_0803_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1605_ ) );
MUX2_X1 \myexu/_4629_ ( .A(\myexu/_2502_ ), .B(\myexu/_1605_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1606_ ) );
AND2_X1 \myexu/_4630_ ( .A1(\myexu/_1606_ ), .A2(\myexu/_0797_ ), .ZN(\myexu/_1607_ ) );
AND2_X2 \myexu/_4631_ ( .A1(\myexu/_0784_ ), .A2(fanout_net_7 ), .ZN(\myexu/_1608_ ) );
NAND2_X1 \myexu/_4632_ ( .A1(\myexu/_1978_ ), .A2(\myexu/_1608_ ), .ZN(\myexu/_1609_ ) );
AND2_X2 \myexu/_4633_ ( .A1(\myexu/_0784_ ), .A2(\myexu/_2118_ ), .ZN(\myexu/_1610_ ) );
INV_X2 \myexu/_4634_ ( .A(\myexu/_1610_ ), .ZN(\myexu/_1611_ ) );
OAI211_X2 \myexu/_4635_ ( .A(\myexu/_1609_ ), .B(\myexu/_2030_ ), .C1(\myexu/_0804_ ), .C2(\myexu/_1611_ ), .ZN(\myexu/_1612_ ) );
OAI221_X1 \myexu/_4636_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2502_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1607_ ), .C2(\myexu/_1612_ ), .ZN(\myexu/_1613_ ) );
OAI21_X1 \myexu/_4637_ ( .A(\myexu/_2303_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1614_ ) );
AOI21_X1 \myexu/_4638_ ( .A(fanout_net_5 ), .B1(\myexu/_1613_ ), .B2(\myexu/_1614_ ), .ZN(\myexu/_0111_ ) );
MUX2_X1 \myexu/_4639_ ( .A(\myexu/_0840_ ), .B(\myexu/_0826_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1615_ ) );
MUX2_X1 \myexu/_4640_ ( .A(\myexu/_2513_ ), .B(\myexu/_1615_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1616_ ) );
AND2_X1 \myexu/_4641_ ( .A1(\myexu/_1616_ ), .A2(\myexu/_0797_ ), .ZN(\myexu/_1617_ ) );
BUF_X4 \myexu/_4642_ ( .A(\myexu/_1608_ ), .Z(\myexu/_1618_ ) );
NAND2_X1 \myexu/_4643_ ( .A1(\myexu/_1995_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1619_ ) );
BUF_X4 \myexu/_4644_ ( .A(\myexu/_1610_ ), .Z(\myexu/_1620_ ) );
NAND2_X1 \myexu/_4645_ ( .A1(\myexu/_0826_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1621_ ) );
NAND3_X1 \myexu/_4646_ ( .A1(\myexu/_1619_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1621_ ), .ZN(\myexu/_1622_ ) );
OAI221_X1 \myexu/_4647_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2513_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1617_ ), .C2(\myexu/_1622_ ), .ZN(\myexu/_1623_ ) );
OAI21_X1 \myexu/_4648_ ( .A(\myexu/_2314_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1624_ ) );
AOI21_X1 \myexu/_4649_ ( .A(fanout_net_5 ), .B1(\myexu/_1623_ ), .B2(\myexu/_1624_ ), .ZN(\myexu/_0112_ ) );
OR2_X1 \myexu/_4650_ ( .A1(\myexu/_1586_ ), .A2(\myexu/_0867_ ), .ZN(\myexu/_1625_ ) );
OAI211_X2 \myexu/_4651_ ( .A(\myexu/_1625_ ), .B(\myexu/_1589_ ), .C1(\myexu/_0852_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1626_ ) );
NAND2_X1 \myexu/_4652_ ( .A1(\myexu/_2516_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1627_ ) );
AOI21_X1 \myexu/_4653_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1626_ ), .B2(\myexu/_1627_ ), .ZN(\myexu/_1628_ ) );
INV_X1 \myexu/_4654_ ( .A(\myexu/_1608_ ), .ZN(\myexu/_1629_ ) );
BUF_X4 \myexu/_4655_ ( .A(\myexu/_1629_ ), .Z(\myexu/_1630_ ) );
OAI221_X1 \myexu/_4656_ ( .A(\myexu/_2030_ ), .B1(\myexu/_0851_ ), .B2(\myexu/_1611_ ), .C1(\myexu/_2011_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1631_ ) );
OAI221_X1 \myexu/_4657_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2516_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1628_ ), .C2(\myexu/_1631_ ), .ZN(\myexu/_1632_ ) );
OAI21_X1 \myexu/_4658_ ( .A(\myexu/_2317_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1633_ ) );
AOI21_X1 \myexu/_4659_ ( .A(fanout_net_5 ), .B1(\myexu/_1632_ ), .B2(\myexu/_1633_ ), .ZN(\myexu/_0113_ ) );
OR2_X1 \myexu/_4660_ ( .A1(\myexu/_1586_ ), .A2(\myexu/_0890_ ), .ZN(\myexu/_1634_ ) );
OAI211_X2 \myexu/_4661_ ( .A(\myexu/_1634_ ), .B(\myexu/_1589_ ), .C1(\myexu/_0875_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1635_ ) );
NAND2_X1 \myexu/_4662_ ( .A1(\myexu/_2517_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1636_ ) );
AOI21_X1 \myexu/_4663_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1635_ ), .B2(\myexu/_1636_ ), .ZN(\myexu/_1637_ ) );
NAND2_X1 \myexu/_4664_ ( .A1(\myexu/_2017_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1638_ ) );
NAND2_X1 \myexu/_4665_ ( .A1(\myexu/_0875_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1639_ ) );
NAND3_X1 \myexu/_4666_ ( .A1(\myexu/_1638_ ), .A2(\myexu/_1639_ ), .A3(\myexu/_2234_ ), .ZN(\myexu/_1640_ ) );
OAI221_X1 \myexu/_4667_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2517_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1637_ ), .C2(\myexu/_1640_ ), .ZN(\myexu/_1641_ ) );
OAI21_X1 \myexu/_4668_ ( .A(\myexu/_2318_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1642_ ) );
AOI21_X1 \myexu/_4669_ ( .A(fanout_net_5 ), .B1(\myexu/_1641_ ), .B2(\myexu/_1642_ ), .ZN(\myexu/_0114_ ) );
BUF_X4 \myexu/_4670_ ( .A(\myexu/_1588_ ), .Z(\myexu/_1643_ ) );
OAI21_X1 \myexu/_4671_ ( .A(\myexu/_0796_ ), .B1(\myexu/_2518_ ), .B2(\myexu/_1643_ ), .ZN(\myexu/_1644_ ) );
MUX2_X1 \myexu/_4672_ ( .A(\myexu/_0909_ ), .B(\myexu/_0904_ ), .S(\myexu/_1586_ ), .Z(\myexu/_1645_ ) );
AOI21_X1 \myexu/_4673_ ( .A(\myexu/_1644_ ), .B1(\myexu/_1645_ ), .B2(\myexu/_1589_ ), .ZN(\myexu/_1646_ ) );
NAND2_X1 \myexu/_4674_ ( .A1(\myexu/_2024_ ), .A2(\myexu/_1608_ ), .ZN(\myexu/_1647_ ) );
OAI211_X2 \myexu/_4675_ ( .A(\myexu/_1647_ ), .B(\myexu/_2030_ ), .C1(\myexu/_0904_ ), .C2(\myexu/_1611_ ), .ZN(\myexu/_1648_ ) );
OAI221_X1 \myexu/_4676_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2518_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1646_ ), .C2(\myexu/_1648_ ), .ZN(\myexu/_1649_ ) );
OAI21_X1 \myexu/_4677_ ( .A(\myexu/_2319_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1650_ ) );
AOI21_X1 \myexu/_4678_ ( .A(fanout_net_6 ), .B1(\myexu/_1649_ ), .B2(\myexu/_1650_ ), .ZN(\myexu/_0115_ ) );
OR2_X1 \myexu/_4679_ ( .A1(\myexu/_1586_ ), .A2(\myexu/_0933_ ), .ZN(\myexu/_1651_ ) );
OAI211_X2 \myexu/_4680_ ( .A(\myexu/_1651_ ), .B(\myexu/_1643_ ), .C1(\myexu/_0926_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1652_ ) );
NAND2_X1 \myexu/_4681_ ( .A1(\myexu/_2519_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1653_ ) );
AOI21_X1 \myexu/_4682_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1652_ ), .B2(\myexu/_1653_ ), .ZN(\myexu/_1654_ ) );
NAND2_X1 \myexu/_4683_ ( .A1(\myexu/_2043_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1655_ ) );
NAND2_X1 \myexu/_4684_ ( .A1(\myexu/_0926_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1656_ ) );
NAND3_X1 \myexu/_4685_ ( .A1(\myexu/_1655_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1656_ ), .ZN(\myexu/_1657_ ) );
OAI221_X1 \myexu/_4686_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2519_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1654_ ), .C2(\myexu/_1657_ ), .ZN(\myexu/_1658_ ) );
OAI21_X1 \myexu/_4687_ ( .A(\myexu/_2320_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1659_ ) );
AOI21_X1 \myexu/_4688_ ( .A(fanout_net_6 ), .B1(\myexu/_1658_ ), .B2(\myexu/_1659_ ), .ZN(\myexu/_0116_ ) );
MUX2_X1 \myexu/_4689_ ( .A(\myexu/_0953_ ), .B(\myexu/_0941_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1660_ ) );
MUX2_X1 \myexu/_4690_ ( .A(\myexu/_2520_ ), .B(\myexu/_1660_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1661_ ) );
AND2_X1 \myexu/_4691_ ( .A1(\myexu/_1661_ ), .A2(\myexu/_0797_ ), .ZN(\myexu/_1662_ ) );
BUF_X4 \myexu/_4692_ ( .A(\myexu/_1610_ ), .Z(\myexu/_1663_ ) );
NAND2_X1 \myexu/_4693_ ( .A1(\myexu/_0941_ ), .A2(\myexu/_1663_ ), .ZN(\myexu/_1664_ ) );
OAI211_X2 \myexu/_4694_ ( .A(\myexu/_2104_ ), .B(\myexu/_1664_ ), .C1(\myexu/_2056_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1665_ ) );
OAI221_X1 \myexu/_4695_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2520_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1662_ ), .C2(\myexu/_1665_ ), .ZN(\myexu/_1666_ ) );
BUF_X4 \myexu/_4696_ ( .A(\myexu/_1598_ ), .Z(\myexu/_1667_ ) );
OAI21_X1 \myexu/_4697_ ( .A(\myexu/_2321_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1668_ ) );
AOI21_X1 \myexu/_4698_ ( .A(fanout_net_6 ), .B1(\myexu/_1666_ ), .B2(\myexu/_1668_ ), .ZN(\myexu/_0117_ ) );
OR2_X1 \myexu/_4699_ ( .A1(\myexu/_1586_ ), .A2(\myexu/_0978_ ), .ZN(\myexu/_1669_ ) );
OAI211_X2 \myexu/_4700_ ( .A(\myexu/_1669_ ), .B(\myexu/_1643_ ), .C1(\myexu/_0971_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1670_ ) );
NAND2_X1 \myexu/_4701_ ( .A1(\myexu/_2521_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1671_ ) );
AOI21_X1 \myexu/_4702_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1670_ ), .B2(\myexu/_1671_ ), .ZN(\myexu/_1672_ ) );
NAND2_X1 \myexu/_4703_ ( .A1(\myexu/_2067_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1673_ ) );
NAND2_X1 \myexu/_4704_ ( .A1(\myexu/_0971_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1674_ ) );
NAND3_X1 \myexu/_4705_ ( .A1(\myexu/_1673_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1674_ ), .ZN(\myexu/_1675_ ) );
OAI221_X1 \myexu/_4706_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2521_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1672_ ), .C2(\myexu/_1675_ ), .ZN(\myexu/_1676_ ) );
BUF_X4 \myexu/_4707_ ( .A(\myexu/_1600_ ), .Z(\myexu/_1677_ ) );
OAI21_X1 \myexu/_4708_ ( .A(\myexu/_2322_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1678_ ) );
AOI21_X1 \myexu/_4709_ ( .A(fanout_net_6 ), .B1(\myexu/_1676_ ), .B2(\myexu/_1678_ ), .ZN(\myexu/_0118_ ) );
OAI21_X1 \myexu/_4710_ ( .A(\myexu/_0796_ ), .B1(\myexu/_2522_ ), .B2(\myexu/_1643_ ), .ZN(\myexu/_1679_ ) );
MUX2_X1 \myexu/_4711_ ( .A(\myexu/_1004_ ), .B(\myexu/_0998_ ), .S(\myexu/_1586_ ), .Z(\myexu/_1680_ ) );
AOI21_X1 \myexu/_4712_ ( .A(\myexu/_1679_ ), .B1(\myexu/_1680_ ), .B2(\myexu/_1589_ ), .ZN(\myexu/_1681_ ) );
OAI221_X1 \myexu/_4713_ ( .A(\myexu/_2030_ ), .B1(\myexu/_0998_ ), .B2(\myexu/_1611_ ), .C1(\myexu/_2079_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1682_ ) );
OAI221_X1 \myexu/_4714_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2522_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1681_ ), .C2(\myexu/_1682_ ), .ZN(\myexu/_1683_ ) );
OAI21_X1 \myexu/_4715_ ( .A(\myexu/_2323_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1684_ ) );
AOI21_X1 \myexu/_4716_ ( .A(fanout_net_6 ), .B1(\myexu/_1683_ ), .B2(\myexu/_1684_ ), .ZN(\myexu/_0119_ ) );
AND2_X1 \myexu/_4717_ ( .A1(\myexu/_1590_ ), .A2(\myexu/_1026_ ), .ZN(\myexu/_1685_ ) );
AOI211_X2 \myexu/_4718_ ( .A(\myexu/_2526_ ), .B(\myexu/_1685_ ), .C1(\myexu/_1019_ ), .C2(\myexu/_1585_ ), .ZN(\myexu/_1686_ ) );
NOR2_X1 \myexu/_4719_ ( .A1(\myexu/_1643_ ), .A2(\myexu/_2492_ ), .ZN(\myexu/_1687_ ) );
NOR3_X1 \myexu/_4720_ ( .A1(\myexu/_1686_ ), .A2(\myexu/_1553_ ), .A3(\myexu/_1687_ ), .ZN(\myexu/_1688_ ) );
NAND3_X1 \myexu/_4721_ ( .A1(\myexu/_2090_ ), .A2(\myexu/_2091_ ), .A3(\myexu/_1618_ ), .ZN(\myexu/_1689_ ) );
NAND2_X1 \myexu/_4722_ ( .A1(\myexu/_1019_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1690_ ) );
NAND3_X1 \myexu/_4723_ ( .A1(\myexu/_1689_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1690_ ), .ZN(\myexu/_1691_ ) );
OAI221_X1 \myexu/_4724_ ( .A(\myexu/_1603_ ), .B1(\myexu/_2492_ ), .B2(\myexu/_1604_ ), .C1(\myexu/_1688_ ), .C2(\myexu/_1691_ ), .ZN(\myexu/_1692_ ) );
OAI21_X1 \myexu/_4725_ ( .A(\myexu/_2293_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1693_ ) );
AOI21_X1 \myexu/_4726_ ( .A(fanout_net_6 ), .B1(\myexu/_1692_ ), .B2(\myexu/_1693_ ), .ZN(\myexu/_0120_ ) );
MUX2_X1 \myexu/_4727_ ( .A(\myexu/_1044_ ), .B(\myexu/_1038_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1694_ ) );
MUX2_X1 \myexu/_4728_ ( .A(\myexu/_2493_ ), .B(\myexu/_1694_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1695_ ) );
AND2_X1 \myexu/_4729_ ( .A1(\myexu/_1695_ ), .A2(\myexu/_0797_ ), .ZN(\myexu/_1696_ ) );
NAND2_X1 \myexu/_4730_ ( .A1(\myexu/_1038_ ), .A2(\myexu/_1663_ ), .ZN(\myexu/_1697_ ) );
OAI211_X2 \myexu/_4731_ ( .A(\myexu/_2104_ ), .B(\myexu/_1697_ ), .C1(\myexu/_2101_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1698_ ) );
OAI221_X1 \myexu/_4732_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2493_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1696_ ), .C2(\myexu/_1698_ ), .ZN(\myexu/_1699_ ) );
OAI21_X1 \myexu/_4733_ ( .A(\myexu/_2294_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1700_ ) );
AOI21_X1 \myexu/_4734_ ( .A(fanout_net_6 ), .B1(\myexu/_1699_ ), .B2(\myexu/_1700_ ), .ZN(\myexu/_0121_ ) );
MUX2_X1 \myexu/_4735_ ( .A(\myexu/_1075_ ), .B(\myexu/_1068_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1701_ ) );
MUX2_X1 \myexu/_4736_ ( .A(\myexu/_2494_ ), .B(\myexu/_1701_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1702_ ) );
AND2_X1 \myexu/_4737_ ( .A1(\myexu/_1702_ ), .A2(\myexu/_0797_ ), .ZN(\myexu/_1703_ ) );
NAND2_X1 \myexu/_4738_ ( .A1(\myexu/_1068_ ), .A2(\myexu/_1663_ ), .ZN(\myexu/_1704_ ) );
OAI211_X2 \myexu/_4739_ ( .A(\myexu/_2104_ ), .B(\myexu/_1704_ ), .C1(\myexu/_0483_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1705_ ) );
OAI221_X1 \myexu/_4740_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2494_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1703_ ), .C2(\myexu/_1705_ ), .ZN(\myexu/_1706_ ) );
OAI21_X1 \myexu/_4741_ ( .A(\myexu/_2295_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1707_ ) );
AOI21_X1 \myexu/_4742_ ( .A(fanout_net_6 ), .B1(\myexu/_1706_ ), .B2(\myexu/_1707_ ), .ZN(\myexu/_0122_ ) );
OR2_X1 \myexu/_4743_ ( .A1(\myexu/_1586_ ), .A2(\myexu/_1096_ ), .ZN(\myexu/_1708_ ) );
OAI211_X2 \myexu/_4744_ ( .A(\myexu/_1708_ ), .B(\myexu/_1643_ ), .C1(\myexu/_1090_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1709_ ) );
NAND2_X1 \myexu/_4745_ ( .A1(\myexu/_2495_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1710_ ) );
AOI21_X1 \myexu/_4746_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1709_ ), .B2(\myexu/_1710_ ), .ZN(\myexu/_1711_ ) );
NAND2_X1 \myexu/_4747_ ( .A1(\myexu/_0491_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1712_ ) );
NAND2_X1 \myexu/_4748_ ( .A1(\myexu/_1090_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1713_ ) );
NAND3_X1 \myexu/_4749_ ( .A1(\myexu/_1712_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1713_ ), .ZN(\myexu/_1714_ ) );
OAI221_X1 \myexu/_4750_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2495_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1711_ ), .C2(\myexu/_1714_ ), .ZN(\myexu/_1715_ ) );
OAI21_X1 \myexu/_4751_ ( .A(\myexu/_2296_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1716_ ) );
AOI21_X1 \myexu/_4752_ ( .A(fanout_net_6 ), .B1(\myexu/_1715_ ), .B2(\myexu/_1716_ ), .ZN(\myexu/_0123_ ) );
MUX2_X1 \myexu/_4753_ ( .A(\myexu/_1119_ ), .B(\myexu/_1110_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1717_ ) );
MUX2_X1 \myexu/_4754_ ( .A(\myexu/_2496_ ), .B(\myexu/_1717_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1718_ ) );
AND2_X1 \myexu/_4755_ ( .A1(\myexu/_1718_ ), .A2(\myexu/_0797_ ), .ZN(\myexu/_1719_ ) );
NAND3_X1 \myexu/_4756_ ( .A1(\myexu/_0498_ ), .A2(\myexu/_0499_ ), .A3(\myexu/_1618_ ), .ZN(\myexu/_1720_ ) );
NAND2_X1 \myexu/_4757_ ( .A1(\myexu/_1110_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1721_ ) );
NAND3_X1 \myexu/_4758_ ( .A1(\myexu/_1720_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1721_ ), .ZN(\myexu/_1722_ ) );
OAI221_X1 \myexu/_4759_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2496_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1719_ ), .C2(\myexu/_1722_ ), .ZN(\myexu/_1723_ ) );
OAI21_X1 \myexu/_4760_ ( .A(\myexu/_2297_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1724_ ) );
AOI21_X1 \myexu/_4761_ ( .A(fanout_net_6 ), .B1(\myexu/_1723_ ), .B2(\myexu/_1724_ ), .ZN(\myexu/_0124_ ) );
AOI21_X1 \myexu/_4762_ ( .A(\myexu/_1267_ ), .B1(\myexu/_2251_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1725_ ) );
MUX2_X1 \myexu/_4763_ ( .A(\myexu/_1138_ ), .B(\myexu/_1132_ ), .S(\myexu/_1585_ ), .Z(\myexu/_1726_ ) );
OAI21_X1 \myexu/_4764_ ( .A(\myexu/_1725_ ), .B1(\myexu/_1726_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1727_ ) );
NOR2_X1 \myexu/_4765_ ( .A1(\myexu/_0505_ ), .A2(\myexu/_1630_ ), .ZN(\myexu/_1728_ ) );
AOI21_X1 \myexu/_4766_ ( .A(\myexu/_1728_ ), .B1(\myexu/_1132_ ), .B2(\myexu/_1620_ ), .ZN(\myexu/_1729_ ) );
NAND3_X1 \myexu/_4767_ ( .A1(\myexu/_1727_ ), .A2(\myexu/_0440_ ), .A3(\myexu/_1729_ ), .ZN(\myexu/_1730_ ) );
OAI211_X2 \myexu/_4768_ ( .A(\myexu/_1730_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2497_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1731_ ) );
OAI21_X1 \myexu/_4769_ ( .A(\myexu/_2298_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1732_ ) );
AOI21_X1 \myexu/_4770_ ( .A(fanout_net_6 ), .B1(\myexu/_1731_ ), .B2(\myexu/_1732_ ), .ZN(\myexu/_0125_ ) );
AND2_X1 \myexu/_4771_ ( .A1(\myexu/_1590_ ), .A2(\myexu/_1173_ ), .ZN(\myexu/_1733_ ) );
AOI211_X2 \myexu/_4772_ ( .A(\myexu/_2526_ ), .B(\myexu/_1733_ ), .C1(\myexu/_1166_ ), .C2(\myexu/_1585_ ), .ZN(\myexu/_1734_ ) );
NOR2_X1 \myexu/_4773_ ( .A1(\myexu/_1643_ ), .A2(\myexu/_2498_ ), .ZN(\myexu/_1735_ ) );
NOR3_X1 \myexu/_4774_ ( .A1(\myexu/_1734_ ), .A2(\myexu/_0787_ ), .A3(\myexu/_1735_ ), .ZN(\myexu/_1736_ ) );
NAND2_X1 \myexu/_4775_ ( .A1(\myexu/_0517_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1737_ ) );
NAND2_X1 \myexu/_4776_ ( .A1(\myexu/_1166_ ), .A2(\myexu/_1620_ ), .ZN(\myexu/_1738_ ) );
NAND3_X1 \myexu/_4777_ ( .A1(\myexu/_1737_ ), .A2(\myexu/_2234_ ), .A3(\myexu/_1738_ ), .ZN(\myexu/_1739_ ) );
OAI221_X1 \myexu/_4778_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2498_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1736_ ), .C2(\myexu/_1739_ ), .ZN(\myexu/_1740_ ) );
OAI21_X1 \myexu/_4779_ ( .A(\myexu/_2299_ ), .B1(\myexu/_1667_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1741_ ) );
AOI21_X1 \myexu/_4780_ ( .A(fanout_net_6 ), .B1(\myexu/_1740_ ), .B2(\myexu/_1741_ ), .ZN(\myexu/_0126_ ) );
NAND2_X1 \myexu/_4781_ ( .A1(\myexu/_1591_ ), .A2(\myexu/_1196_ ), .ZN(\myexu/_1742_ ) );
OAI211_X2 \myexu/_4782_ ( .A(\myexu/_1742_ ), .B(\myexu/_1643_ ), .C1(\myexu/_1190_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1743_ ) );
NAND2_X1 \myexu/_4783_ ( .A1(\myexu/_2499_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1744_ ) );
AOI21_X1 \myexu/_4784_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1743_ ), .B2(\myexu/_1744_ ), .ZN(\myexu/_1745_ ) );
NAND2_X1 \myexu/_4785_ ( .A1(\myexu/_1190_ ), .A2(\myexu/_1663_ ), .ZN(\myexu/_1746_ ) );
OAI211_X2 \myexu/_4786_ ( .A(\myexu/_2104_ ), .B(\myexu/_1746_ ), .C1(\myexu/_0526_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1747_ ) );
OAI221_X1 \myexu/_4787_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2499_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1745_ ), .C2(\myexu/_1747_ ), .ZN(\myexu/_1748_ ) );
BUF_X4 \myexu/_4788_ ( .A(\myexu/_1598_ ), .Z(\myexu/_1749_ ) );
OAI21_X1 \myexu/_4789_ ( .A(\myexu/_2300_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1677_ ), .ZN(\myexu/_1750_ ) );
AOI21_X1 \myexu/_4790_ ( .A(fanout_net_6 ), .B1(\myexu/_1748_ ), .B2(\myexu/_1750_ ), .ZN(\myexu/_0127_ ) );
AOI221_X4 \myexu/_4791_ ( .A(\myexu/_2028_ ), .B1(\myexu/_1215_ ), .B2(\myexu/_1610_ ), .C1(\myexu/_0535_ ), .C2(\myexu/_1608_ ), .ZN(\myexu/_1751_ ) );
AND2_X1 \myexu/_4792_ ( .A1(\myexu/_1590_ ), .A2(\myexu/_1222_ ), .ZN(\myexu/_1752_ ) );
AOI211_X2 \myexu/_4793_ ( .A(\myexu/_2526_ ), .B(\myexu/_1752_ ), .C1(\myexu/_1215_ ), .C2(\myexu/_1585_ ), .ZN(\myexu/_1753_ ) );
OAI21_X1 \myexu/_4794_ ( .A(\myexu/_0796_ ), .B1(\myexu/_2500_ ), .B2(\myexu/_1643_ ), .ZN(\myexu/_1754_ ) );
OAI21_X1 \myexu/_4795_ ( .A(\myexu/_1751_ ), .B1(\myexu/_1753_ ), .B2(\myexu/_1754_ ), .ZN(\myexu/_1755_ ) );
OAI211_X2 \myexu/_4796_ ( .A(\myexu/_1755_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2500_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1756_ ) );
BUF_X4 \myexu/_4797_ ( .A(\myexu/_1600_ ), .Z(\myexu/_1757_ ) );
OAI21_X1 \myexu/_4798_ ( .A(\myexu/_2301_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1758_ ) );
AOI21_X1 \myexu/_4799_ ( .A(fanout_net_6 ), .B1(\myexu/_1756_ ), .B2(\myexu/_1758_ ), .ZN(\myexu/_0128_ ) );
AOI21_X1 \myexu/_4800_ ( .A(\myexu/_1267_ ), .B1(\myexu/_0349_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1759_ ) );
MUX2_X1 \myexu/_4801_ ( .A(\myexu/_1242_ ), .B(\myexu/_1236_ ), .S(\myexu/_1585_ ), .Z(\myexu/_1760_ ) );
OAI21_X1 \myexu/_4802_ ( .A(\myexu/_1759_ ), .B1(\myexu/_1760_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1761_ ) );
NOR2_X1 \myexu/_4803_ ( .A1(\myexu/_0542_ ), .A2(\myexu/_1630_ ), .ZN(\myexu/_1762_ ) );
AOI21_X1 \myexu/_4804_ ( .A(\myexu/_1762_ ), .B1(\myexu/_1236_ ), .B2(\myexu/_1620_ ), .ZN(\myexu/_1763_ ) );
NAND3_X1 \myexu/_4805_ ( .A1(\myexu/_1761_ ), .A2(\myexu/_0440_ ), .A3(\myexu/_1763_ ), .ZN(\myexu/_1764_ ) );
OAI211_X2 \myexu/_4806_ ( .A(\myexu/_1764_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2501_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1765_ ) );
OAI21_X1 \myexu/_4807_ ( .A(\myexu/_2302_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1766_ ) );
AOI21_X1 \myexu/_4808_ ( .A(fanout_net_6 ), .B1(\myexu/_1765_ ), .B2(\myexu/_1766_ ), .ZN(\myexu/_0129_ ) );
NAND2_X1 \myexu/_4809_ ( .A1(\myexu/_1590_ ), .A2(\myexu/_1270_ ), .ZN(\myexu/_1767_ ) );
OAI211_X2 \myexu/_4810_ ( .A(\myexu/_1767_ ), .B(\myexu/_1643_ ), .C1(\myexu/_1262_ ), .C2(\myexu/_1591_ ), .ZN(\myexu/_1768_ ) );
NAND2_X1 \myexu/_4811_ ( .A1(\myexu/_2503_ ), .A2(\myexu/_2526_ ), .ZN(\myexu/_1769_ ) );
AOI21_X1 \myexu/_4812_ ( .A(\myexu/_1553_ ), .B1(\myexu/_1768_ ), .B2(\myexu/_1769_ ), .ZN(\myexu/_1770_ ) );
NAND2_X1 \myexu/_4813_ ( .A1(\myexu/_1262_ ), .A2(\myexu/_1663_ ), .ZN(\myexu/_1771_ ) );
OAI211_X2 \myexu/_4814_ ( .A(\myexu/_2104_ ), .B(\myexu/_1771_ ), .C1(\myexu/_0555_ ), .C2(\myexu/_1630_ ), .ZN(\myexu/_1772_ ) );
OAI221_X1 \myexu/_4815_ ( .A(\myexu/_1550_ ), .B1(\myexu/_2503_ ), .B2(\myexu/_2031_ ), .C1(\myexu/_1770_ ), .C2(\myexu/_1772_ ), .ZN(\myexu/_1773_ ) );
OAI21_X1 \myexu/_4816_ ( .A(\myexu/_2304_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1774_ ) );
AOI21_X1 \myexu/_4817_ ( .A(fanout_net_6 ), .B1(\myexu/_1773_ ), .B2(\myexu/_1774_ ), .ZN(\myexu/_0130_ ) );
AOI21_X1 \myexu/_4818_ ( .A(\myexu/_1267_ ), .B1(\myexu/_0368_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1775_ ) );
MUX2_X1 \myexu/_4819_ ( .A(\myexu/_1275_ ), .B(\myexu/_1291_ ), .S(\myexu/_1585_ ), .Z(\myexu/_1776_ ) );
OAI21_X1 \myexu/_4820_ ( .A(\myexu/_1775_ ), .B1(\myexu/_1776_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1777_ ) );
NOR2_X1 \myexu/_4821_ ( .A1(\myexu/_0561_ ), .A2(\myexu/_1630_ ), .ZN(\myexu/_1778_ ) );
AOI21_X1 \myexu/_4822_ ( .A(\myexu/_1778_ ), .B1(\myexu/_1291_ ), .B2(\myexu/_1663_ ), .ZN(\myexu/_1779_ ) );
NAND3_X1 \myexu/_4823_ ( .A1(\myexu/_1777_ ), .A2(\myexu/_0440_ ), .A3(\myexu/_1779_ ), .ZN(\myexu/_1780_ ) );
OAI211_X2 \myexu/_4824_ ( .A(\myexu/_1780_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2504_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1781_ ) );
OAI21_X1 \myexu/_4825_ ( .A(\myexu/_2305_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1782_ ) );
AOI21_X1 \myexu/_4826_ ( .A(fanout_net_6 ), .B1(\myexu/_1781_ ), .B2(\myexu/_1782_ ), .ZN(\myexu/_0131_ ) );
AOI21_X1 \myexu/_4827_ ( .A(\myexu/_1267_ ), .B1(\myexu/_1300_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1783_ ) );
MUX2_X1 \myexu/_4828_ ( .A(\myexu/_1322_ ), .B(\myexu/_1314_ ), .S(\myexu/_1585_ ), .Z(\myexu/_1784_ ) );
OAI21_X1 \myexu/_4829_ ( .A(\myexu/_1783_ ), .B1(\myexu/_1784_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1785_ ) );
NOR2_X1 \myexu/_4830_ ( .A1(\myexu/_0569_ ), .A2(\myexu/_1629_ ), .ZN(\myexu/_1786_ ) );
AOI21_X1 \myexu/_4831_ ( .A(\myexu/_1786_ ), .B1(\myexu/_1314_ ), .B2(\myexu/_1663_ ), .ZN(\myexu/_1787_ ) );
NAND3_X1 \myexu/_4832_ ( .A1(\myexu/_1785_ ), .A2(\myexu/_0440_ ), .A3(\myexu/_1787_ ), .ZN(\myexu/_1788_ ) );
OAI211_X2 \myexu/_4833_ ( .A(\myexu/_1788_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2505_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1789_ ) );
OAI21_X1 \myexu/_4834_ ( .A(\myexu/_2306_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1790_ ) );
AOI21_X1 \myexu/_4835_ ( .A(fanout_net_6 ), .B1(\myexu/_1789_ ), .B2(\myexu/_1790_ ), .ZN(\myexu/_0132_ ) );
OAI21_X1 \myexu/_4836_ ( .A(\myexu/_0785_ ), .B1(\myexu/_1336_ ), .B2(fanout_net_7 ), .ZN(\myexu/_1791_ ) );
AOI21_X1 \myexu/_4837_ ( .A(\myexu/_1791_ ), .B1(\myexu/_0575_ ), .B2(fanout_net_7 ), .ZN(\myexu/_1792_ ) );
MUX2_X1 \myexu/_4838_ ( .A(\myexu/_1342_ ), .B(\myexu/_1336_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1793_ ) );
MUX2_X2 \myexu/_4839_ ( .A(\myexu/_2506_ ), .B(\myexu/_1793_ ), .S(\myexu/_0762_ ), .Z(\myexu/_1794_ ) );
AOI21_X1 \myexu/_4840_ ( .A(\myexu/_1792_ ), .B1(\myexu/_1794_ ), .B2(\myexu/_0795_ ), .ZN(\myexu/_1795_ ) );
MUX2_X2 \myexu/_4841_ ( .A(\myexu/_0385_ ), .B(\myexu/_1795_ ), .S(\myexu/_2029_ ), .Z(\myexu/_1796_ ) );
OR3_X2 \myexu/_4842_ ( .A1(\myexu/_1796_ ), .A2(\myexu/_1600_ ), .A3(\myexu/_1598_ ), .ZN(\myexu/_1797_ ) );
OAI21_X1 \myexu/_4843_ ( .A(\myexu/_2307_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1798_ ) );
AOI21_X1 \myexu/_4844_ ( .A(fanout_net_6 ), .B1(\myexu/_1797_ ), .B2(\myexu/_1798_ ), .ZN(\myexu/_0133_ ) );
OAI21_X1 \myexu/_4845_ ( .A(\myexu/_0795_ ), .B1(\myexu/_2507_ ), .B2(\myexu/_0762_ ), .ZN(\myexu/_1799_ ) );
OAI21_X1 \myexu/_4846_ ( .A(\myexu/_1611_ ), .B1(\myexu/_1590_ ), .B2(\myexu/_1799_ ), .ZN(\myexu/_1800_ ) );
AOI221_X2 \myexu/_4847_ ( .A(\myexu/_2028_ ), .B1(\myexu/_0588_ ), .B2(\myexu/_1608_ ), .C1(\myexu/_1800_ ), .C2(\myexu/_1367_ ), .ZN(\myexu/_1801_ ) );
AOI21_X1 \myexu/_4848_ ( .A(\myexu/_2526_ ), .B1(\myexu/_1591_ ), .B2(\myexu/_1374_ ), .ZN(\myexu/_1802_ ) );
OAI21_X1 \myexu/_4849_ ( .A(\myexu/_1801_ ), .B1(\myexu/_1799_ ), .B2(\myexu/_1802_ ), .ZN(\myexu/_1803_ ) );
OAI211_X2 \myexu/_4850_ ( .A(\myexu/_1803_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2507_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1804_ ) );
OAI21_X1 \myexu/_4851_ ( .A(\myexu/_2308_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1805_ ) );
AOI21_X1 \myexu/_4852_ ( .A(fanout_net_6 ), .B1(\myexu/_1804_ ), .B2(\myexu/_1805_ ), .ZN(\myexu/_0134_ ) );
OAI21_X1 \myexu/_4853_ ( .A(\myexu/_0785_ ), .B1(\myexu/_1394_ ), .B2(fanout_net_7 ), .ZN(\myexu/_1806_ ) );
AOI21_X1 \myexu/_4854_ ( .A(\myexu/_1806_ ), .B1(\myexu/_0594_ ), .B2(\myexu/_2523_ ), .ZN(\myexu/_1807_ ) );
MUX2_X1 \myexu/_4855_ ( .A(\myexu/_1401_ ), .B(\myexu/_1394_ ), .S(\myexu/_1584_ ), .Z(\myexu/_1808_ ) );
MUX2_X2 \myexu/_4856_ ( .A(\myexu/_2508_ ), .B(\myexu/_1808_ ), .S(\myexu/_0762_ ), .Z(\myexu/_1809_ ) );
AOI21_X1 \myexu/_4857_ ( .A(\myexu/_1807_ ), .B1(\myexu/_1809_ ), .B2(\myexu/_0795_ ), .ZN(\myexu/_1810_ ) );
MUX2_X2 \myexu/_4858_ ( .A(\myexu/_0401_ ), .B(\myexu/_1810_ ), .S(\myexu/_2029_ ), .Z(\myexu/_1811_ ) );
OR3_X2 \myexu/_4859_ ( .A1(\myexu/_1811_ ), .A2(\myexu/_1600_ ), .A3(\myexu/_1598_ ), .ZN(\myexu/_1812_ ) );
OAI21_X1 \myexu/_4860_ ( .A(\myexu/_2309_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1813_ ) );
AOI21_X1 \myexu/_4861_ ( .A(fanout_net_6 ), .B1(\myexu/_1812_ ), .B2(\myexu/_1813_ ), .ZN(\myexu/_0135_ ) );
AOI21_X1 \myexu/_4862_ ( .A(\myexu/_0786_ ), .B1(\myexu/_0411_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1814_ ) );
MUX2_X1 \myexu/_4863_ ( .A(\myexu/_1424_ ), .B(\myexu/_1416_ ), .S(\myexu/_1585_ ), .Z(\myexu/_1815_ ) );
OAI21_X1 \myexu/_4864_ ( .A(\myexu/_1814_ ), .B1(\myexu/_1815_ ), .B2(\myexu/_2526_ ), .ZN(\myexu/_1816_ ) );
NOR2_X1 \myexu/_4865_ ( .A1(\myexu/_0601_ ), .A2(\myexu/_1629_ ), .ZN(\myexu/_1817_ ) );
AOI21_X1 \myexu/_4866_ ( .A(\myexu/_1817_ ), .B1(\myexu/_1416_ ), .B2(\myexu/_1663_ ), .ZN(\myexu/_1818_ ) );
NAND3_X1 \myexu/_4867_ ( .A1(\myexu/_1816_ ), .A2(\myexu/_0440_ ), .A3(\myexu/_1818_ ), .ZN(\myexu/_1819_ ) );
OAI211_X2 \myexu/_4868_ ( .A(\myexu/_1819_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2509_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1820_ ) );
OAI21_X1 \myexu/_4869_ ( .A(\myexu/_2310_ ), .B1(\myexu/_1749_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1821_ ) );
AOI21_X1 \myexu/_4870_ ( .A(fanout_net_6 ), .B1(\myexu/_1820_ ), .B2(\myexu/_1821_ ), .ZN(\myexu/_0136_ ) );
OAI21_X1 \myexu/_4871_ ( .A(\myexu/_0784_ ), .B1(\myexu/_1438_ ), .B2(\myexu/_2523_ ), .ZN(\myexu/_1822_ ) );
AOI21_X1 \myexu/_4872_ ( .A(\myexu/_1822_ ), .B1(\myexu/_0607_ ), .B2(\myexu/_2523_ ), .ZN(\myexu/_1823_ ) );
MUX2_X1 \myexu/_4873_ ( .A(\myexu/_1444_ ), .B(\myexu/_1438_ ), .S(\myexu/_1583_ ), .Z(\myexu/_1824_ ) );
MUX2_X1 \myexu/_4874_ ( .A(\myexu/_2510_ ), .B(\myexu/_1824_ ), .S(\myexu/_0762_ ), .Z(\myexu/_1825_ ) );
AOI21_X1 \myexu/_4875_ ( .A(\myexu/_1823_ ), .B1(\myexu/_1825_ ), .B2(\myexu/_0795_ ), .ZN(\myexu/_1826_ ) );
MUX2_X1 \myexu/_4876_ ( .A(\myexu/_1447_ ), .B(\myexu/_1826_ ), .S(\myexu/_2029_ ), .Z(\myexu/_1827_ ) );
OR3_X1 \myexu/_4877_ ( .A1(\myexu/_1827_ ), .A2(\myexu/_1600_ ), .A3(\myexu/_1598_ ), .ZN(\myexu/_1828_ ) );
OAI21_X1 \myexu/_4878_ ( .A(\myexu/_2311_ ), .B1(\myexu/_1598_ ), .B2(\myexu/_1757_ ), .ZN(\myexu/_1829_ ) );
AOI21_X1 \myexu/_4879_ ( .A(fanout_net_6 ), .B1(\myexu/_1828_ ), .B2(\myexu/_1829_ ), .ZN(\myexu/_0137_ ) );
NOR4_X1 \myexu/_4880_ ( .A1(\myexu/_1963_ ), .A2(\myexu/_0816_ ), .A3(\myexu/_0637_ ), .A4(\myexu/_2511_ ), .ZN(\myexu/_1830_ ) );
NOR3_X1 \myexu/_4881_ ( .A1(\myexu/_1830_ ), .A2(\myexu/_1600_ ), .A3(\myexu/_1598_ ), .ZN(\myexu/_1831_ ) );
OAI21_X1 \myexu/_4882_ ( .A(\myexu/_0797_ ), .B1(\myexu/_2511_ ), .B2(\myexu/_1589_ ), .ZN(\myexu/_1832_ ) );
MUX2_X1 \myexu/_4883_ ( .A(\myexu/_1471_ ), .B(\myexu/_1465_ ), .S(\myexu/_1586_ ), .Z(\myexu/_1833_ ) );
AOI21_X1 \myexu/_4884_ ( .A(\myexu/_1832_ ), .B1(\myexu/_1833_ ), .B2(\myexu/_1589_ ), .ZN(\myexu/_1834_ ) );
NAND2_X1 \myexu/_4885_ ( .A1(\myexu/_0614_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1835_ ) );
OAI211_X2 \myexu/_4886_ ( .A(\myexu/_1835_ ), .B(\myexu/_0440_ ), .C1(\myexu/_1465_ ), .C2(\myexu/_1611_ ), .ZN(\myexu/_1836_ ) );
OAI21_X1 \myexu/_4887_ ( .A(\myexu/_1831_ ), .B1(\myexu/_1834_ ), .B2(\myexu/_1836_ ), .ZN(\myexu/_1837_ ) );
CLKBUF_X2 \myexu/_4888_ ( .A(\myexu/_1972_ ), .Z(\myexu/_1838_ ) );
OAI21_X1 \myexu/_4889_ ( .A(\myexu/_2312_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1839_ ) );
NAND3_X1 \myexu/_4890_ ( .A1(\myexu/_1837_ ), .A2(\myexu/_1838_ ), .A3(\myexu/_1839_ ), .ZN(\myexu/_0138_ ) );
AOI211_X4 \myexu/_4891_ ( .A(\myexu/_1600_ ), .B(\myexu/_1548_ ), .C1(\myexu/_0449_ ), .C2(\myexu/_2133_ ), .ZN(\myexu/_1840_ ) );
OAI21_X1 \myexu/_4892_ ( .A(\myexu/_0797_ ), .B1(\myexu/_2512_ ), .B2(\myexu/_1589_ ), .ZN(\myexu/_1841_ ) );
INV_X1 \myexu/_4893_ ( .A(\myexu/_1486_ ), .ZN(\myexu/_1842_ ) );
MUX2_X1 \myexu/_4894_ ( .A(\myexu/_1493_ ), .B(\myexu/_1842_ ), .S(\myexu/_1586_ ), .Z(\myexu/_1843_ ) );
AOI21_X1 \myexu/_4895_ ( .A(\myexu/_1841_ ), .B1(\myexu/_1843_ ), .B2(\myexu/_1589_ ), .ZN(\myexu/_1844_ ) );
NAND2_X1 \myexu/_4896_ ( .A1(\myexu/_0621_ ), .A2(\myexu/_1618_ ), .ZN(\myexu/_1845_ ) );
OAI211_X2 \myexu/_4897_ ( .A(\myexu/_1845_ ), .B(\myexu/_0440_ ), .C1(\myexu/_1842_ ), .C2(\myexu/_1611_ ), .ZN(\myexu/_1846_ ) );
OAI21_X1 \myexu/_4898_ ( .A(\myexu/_1840_ ), .B1(\myexu/_1844_ ), .B2(\myexu/_1846_ ), .ZN(\myexu/_1847_ ) );
OAI21_X1 \myexu/_4899_ ( .A(\myexu/_2313_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1601_ ), .ZN(\myexu/_1848_ ) );
NAND3_X1 \myexu/_4900_ ( .A1(\myexu/_1847_ ), .A2(\myexu/_1838_ ), .A3(\myexu/_1848_ ), .ZN(\myexu/_0139_ ) );
AOI22_X1 \myexu/_4901_ ( .A1(\myexu/_0627_ ), .A2(\myexu/_1608_ ), .B1(\myexu/_1522_ ), .B2(\myexu/_1663_ ), .ZN(\myexu/_1849_ ) );
AND2_X2 \myexu/_4902_ ( .A1(\myexu/_1590_ ), .A2(\myexu/_1506_ ), .ZN(\myexu/_1850_ ) );
AOI211_X2 \myexu/_4903_ ( .A(\myexu/_2526_ ), .B(\myexu/_1850_ ), .C1(\myexu/_1522_ ), .C2(\myexu/_1585_ ), .ZN(\myexu/_1851_ ) );
OAI21_X1 \myexu/_4904_ ( .A(\myexu/_0796_ ), .B1(\myexu/_2514_ ), .B2(\myexu/_1588_ ), .ZN(\myexu/_1852_ ) );
OAI211_X2 \myexu/_4905_ ( .A(\myexu/_0440_ ), .B(\myexu/_1849_ ), .C1(\myexu/_1851_ ), .C2(\myexu/_1852_ ), .ZN(\myexu/_1853_ ) );
OAI211_X2 \myexu/_4906_ ( .A(\myexu/_1853_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2514_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1854_ ) );
OAI21_X1 \myexu/_4907_ ( .A(\myexu/_2315_ ), .B1(\myexu/_1598_ ), .B2(\myexu/_1600_ ), .ZN(\myexu/_1855_ ) );
AOI21_X1 \myexu/_4908_ ( .A(fanout_net_6 ), .B1(\myexu/_1854_ ), .B2(\myexu/_1855_ ), .ZN(\myexu/_0140_ ) );
NOR2_X1 \myexu/_4909_ ( .A1(\myexu/_0633_ ), .A2(\myexu/_1629_ ), .ZN(\myexu/_1856_ ) );
AOI21_X1 \myexu/_4910_ ( .A(\myexu/_1856_ ), .B1(\myexu/_1538_ ), .B2(\myexu/_1663_ ), .ZN(\myexu/_1857_ ) );
NAND2_X1 \myexu/_4911_ ( .A1(\myexu/_1590_ ), .A2(\myexu/_1545_ ), .ZN(\myexu/_1858_ ) );
OAI21_X1 \myexu/_4912_ ( .A(\myexu/_1858_ ), .B1(\myexu/_1538_ ), .B2(\myexu/_1590_ ), .ZN(\myexu/_1859_ ) );
MUX2_X2 \myexu/_4913_ ( .A(\myexu/_0466_ ), .B(\myexu/_1859_ ), .S(\myexu/_1588_ ), .Z(\myexu/_1860_ ) );
OAI211_X2 \myexu/_4914_ ( .A(\myexu/_2234_ ), .B(\myexu/_1857_ ), .C1(\myexu/_1860_ ), .C2(\myexu/_1553_ ), .ZN(\myexu/_1861_ ) );
OAI211_X2 \myexu/_4915_ ( .A(\myexu/_1861_ ), .B(\myexu/_1551_ ), .C1(\myexu/_2515_ ), .C2(\myexu/_1552_ ), .ZN(\myexu/_1862_ ) );
OAI21_X1 \myexu/_4916_ ( .A(\myexu/_2316_ ), .B1(\myexu/_1598_ ), .B2(\myexu/_1600_ ), .ZN(\myexu/_1863_ ) );
AOI21_X1 \myexu/_4917_ ( .A(fanout_net_6 ), .B1(\myexu/_1862_ ), .B2(\myexu/_1863_ ), .ZN(\myexu/_0141_ ) );
INV_X1 \myexu/_4918_ ( .A(\myexu/_0242_ ), .ZN(\myexu/_1864_ ) );
OR2_X1 \myexu/_4919_ ( .A1(\myexu/_1864_ ), .A2(\myexu/_0241_ ), .ZN(\myexu/_1865_ ) );
AOI221_X4 \myexu/_4920_ ( .A(\myexu/_1982_ ), .B1(\myexu/_2528_ ), .B2(\myexu/_1958_ ), .C1(\myexu/_0786_ ), .C2(\myexu/_2523_ ), .ZN(\myexu/_1866_ ) );
OAI22_X1 \myexu/_4921_ ( .A1(\myexu/_2529_ ), .A2(\myexu/_0637_ ), .B1(\myexu/_1864_ ), .B2(\myexu/_0241_ ), .ZN(\myexu/_1867_ ) );
OAI211_X2 \myexu/_4922_ ( .A(\myexu/_0816_ ), .B(\myexu/_2530_ ), .C1(\myexu/_2527_ ), .C2(\myexu/_2528_ ), .ZN(\myexu/_1868_ ) );
NAND2_X1 \myexu/_4923_ ( .A1(\myexu/_1867_ ), .A2(\myexu/_1868_ ), .ZN(\myexu/_1869_ ) );
AOI221_X4 \myexu/_4924_ ( .A(fanout_net_6 ), .B1(\myexu/_1982_ ), .B2(\myexu/_1865_ ), .C1(\myexu/_1866_ ), .C2(\myexu/_1869_ ), .ZN(\myexu/_0142_ ) );
BUF_X4 \myexu/_4925_ ( .A(\myexu/_1981_ ), .Z(\myexu/_1870_ ) );
NOR2_X1 \myexu/_4926_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2324_ ), .ZN(\myexu/_1871_ ) );
AOI211_X4 \myexu/_4927_ ( .A(fanout_net_6 ), .B(\myexu/_1871_ ), .C1(\myexu/_2105_ ), .C2(\myexu/_2003_ ), .ZN(\myexu/_0143_ ) );
MUX2_X1 \myexu/_4928_ ( .A(\myexu/_2335_ ), .B(\myexu/_2271_ ), .S(\myexu/_1987_ ), .Z(\myexu/_1872_ ) );
AND2_X1 \myexu/_4929_ ( .A1(\myexu/_1872_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0144_ ) );
NOR2_X1 \myexu/_4930_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2346_ ), .ZN(\myexu/_1873_ ) );
AOI211_X4 \myexu/_4931_ ( .A(fanout_net_6 ), .B(\myexu/_1873_ ), .C1(\myexu/_0840_ ), .C2(\myexu/_2003_ ), .ZN(\myexu/_0145_ ) );
NOR2_X1 \myexu/_4932_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2349_ ), .ZN(\myexu/_1874_ ) );
AOI211_X4 \myexu/_4933_ ( .A(fanout_net_6 ), .B(\myexu/_1874_ ), .C1(\myexu/_2150_ ), .C2(\myexu/_2003_ ), .ZN(\myexu/_0146_ ) );
NOR2_X1 \myexu/_4934_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2350_ ), .ZN(\myexu/_1875_ ) );
AOI211_X4 \myexu/_4935_ ( .A(fanout_net_6 ), .B(\myexu/_1875_ ), .C1(\myexu/_0889_ ), .C2(\myexu/_2003_ ), .ZN(\myexu/_0147_ ) );
MUX2_X1 \myexu/_4936_ ( .A(\myexu/_2351_ ), .B(\myexu/_2287_ ), .S(\myexu/_1987_ ), .Z(\myexu/_1876_ ) );
AND2_X1 \myexu/_4937_ ( .A1(\myexu/_1876_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0148_ ) );
NOR2_X1 \myexu/_4938_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2352_ ), .ZN(\myexu/_1877_ ) );
AOI211_X4 \myexu/_4939_ ( .A(\myexu/_2426_ ), .B(\myexu/_1877_ ), .C1(\myexu/_2177_ ), .C2(\myexu/_2003_ ), .ZN(\myexu/_0149_ ) );
NOR2_X1 \myexu/_4940_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2353_ ), .ZN(\myexu/_1878_ ) );
BUF_X4 \myexu/_4941_ ( .A(\myexu/_1981_ ), .Z(\myexu/_1879_ ) );
AOI211_X4 \myexu/_4942_ ( .A(\myexu/_2426_ ), .B(\myexu/_1878_ ), .C1(\myexu/_0952_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0150_ ) );
NOR2_X1 \myexu/_4943_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2354_ ), .ZN(\myexu/_1880_ ) );
AOI211_X4 \myexu/_4944_ ( .A(\myexu/_2426_ ), .B(\myexu/_1880_ ), .C1(\myexu/_0977_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0151_ ) );
NOR2_X1 \myexu/_4945_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2355_ ), .ZN(\myexu/_1881_ ) );
AOI211_X4 \myexu/_4946_ ( .A(\myexu/_2426_ ), .B(\myexu/_1881_ ), .C1(\myexu/_2203_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0152_ ) );
NOR2_X1 \myexu/_4947_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2325_ ), .ZN(\myexu/_1882_ ) );
AOI211_X4 \myexu/_4948_ ( .A(\myexu/_2426_ ), .B(\myexu/_1882_ ), .C1(\myexu/_1025_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0153_ ) );
MUX2_X1 \myexu/_4949_ ( .A(\myexu/_2326_ ), .B(\myexu/_2262_ ), .S(\myexu/_1987_ ), .Z(\myexu/_1883_ ) );
AND2_X1 \myexu/_4950_ ( .A1(\myexu/_1883_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0154_ ) );
NOR2_X1 \myexu/_4951_ ( .A1(\myexu/_1870_ ), .A2(\myexu/_2327_ ), .ZN(\myexu/_1884_ ) );
AOI211_X4 \myexu/_4952_ ( .A(\myexu/_2426_ ), .B(\myexu/_1884_ ), .C1(\myexu/_1074_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0155_ ) );
BUF_X4 \myexu/_4953_ ( .A(\myexu/_1981_ ), .Z(\myexu/_1885_ ) );
NOR2_X1 \myexu/_4954_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2328_ ), .ZN(\myexu/_1886_ ) );
AOI211_X4 \myexu/_4955_ ( .A(\myexu/_2426_ ), .B(\myexu/_1886_ ), .C1(\myexu/_2233_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0156_ ) );
NOR2_X1 \myexu/_4956_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2329_ ), .ZN(\myexu/_1887_ ) );
AOI211_X4 \myexu/_4957_ ( .A(\myexu/_2426_ ), .B(\myexu/_1887_ ), .C1(\myexu/_1118_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0157_ ) );
NOR2_X1 \myexu/_4958_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2330_ ), .ZN(\myexu/_1888_ ) );
AOI211_X4 \myexu/_4959_ ( .A(\myexu/_2426_ ), .B(\myexu/_1888_ ), .C1(\myexu/_2256_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0158_ ) );
NOR2_X1 \myexu/_4960_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2331_ ), .ZN(\myexu/_1889_ ) );
AOI211_X4 \myexu/_4961_ ( .A(\myexu/_2426_ ), .B(\myexu/_1889_ ), .C1(\myexu/_1194_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0159_ ) );
MUX2_X1 \myexu/_4962_ ( .A(\myexu/_2332_ ), .B(\myexu/_2268_ ), .S(\myexu/_1987_ ), .Z(\myexu/_1890_ ) );
AND2_X1 \myexu/_4963_ ( .A1(\myexu/_1890_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0160_ ) );
BUF_X4 \myexu/_4964_ ( .A(\myexu/_1981_ ), .Z(\myexu/_1891_ ) );
MUX2_X1 \myexu/_4965_ ( .A(\myexu/_2333_ ), .B(\myexu/_2269_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1892_ ) );
AND2_X1 \myexu/_4966_ ( .A1(\myexu/_1892_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0161_ ) );
NOR2_X1 \myexu/_4967_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2334_ ), .ZN(\myexu/_1893_ ) );
AOI211_X4 \myexu/_4968_ ( .A(\myexu/_2426_ ), .B(\myexu/_1893_ ), .C1(\myexu/_0354_ ), .C2(\myexu/_1879_ ), .ZN(\myexu/_0162_ ) );
NOR2_X1 \myexu/_4969_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2336_ ), .ZN(\myexu/_1894_ ) );
BUF_X4 \myexu/_4970_ ( .A(\myexu/_1981_ ), .Z(\myexu/_1895_ ) );
AOI211_X4 \myexu/_4971_ ( .A(\myexu/_2426_ ), .B(\myexu/_1894_ ), .C1(\myexu/_1273_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0163_ ) );
NOR2_X1 \myexu/_4972_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2337_ ), .ZN(\myexu/_1896_ ) );
AOI211_X4 \myexu/_4973_ ( .A(\myexu/_2426_ ), .B(\myexu/_1896_ ), .C1(\myexu/_0364_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0164_ ) );
MUX2_X1 \myexu/_4974_ ( .A(\myexu/_2338_ ), .B(\myexu/_2274_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1897_ ) );
AND2_X1 \myexu/_4975_ ( .A1(\myexu/_1897_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0165_ ) );
MUX2_X1 \myexu/_4976_ ( .A(\myexu/_2339_ ), .B(\myexu/_2275_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1898_ ) );
AND2_X1 \myexu/_4977_ ( .A1(\myexu/_1898_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0166_ ) );
NOR2_X1 \myexu/_4978_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2340_ ), .ZN(\myexu/_1899_ ) );
AOI211_X4 \myexu/_4979_ ( .A(\myexu/_2426_ ), .B(\myexu/_1899_ ), .C1(\myexu/_1399_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0167_ ) );
NOR2_X1 \myexu/_4980_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2341_ ), .ZN(\myexu/_1900_ ) );
AOI211_X4 \myexu/_4981_ ( .A(\myexu/_2426_ ), .B(\myexu/_1900_ ), .C1(\myexu/_0406_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0168_ ) );
NOR2_X1 \myexu/_4982_ ( .A1(\myexu/_1885_ ), .A2(\myexu/_2342_ ), .ZN(\myexu/_1901_ ) );
AOI211_X4 \myexu/_4983_ ( .A(\myexu/_2426_ ), .B(\myexu/_1901_ ), .C1(\myexu/_1423_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0169_ ) );
NOR2_X1 \myexu/_4984_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2343_ ), .ZN(\myexu/_1902_ ) );
AOI211_X4 \myexu/_4985_ ( .A(\myexu/_2426_ ), .B(\myexu/_1902_ ), .C1(\myexu/_0419_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0170_ ) );
MUX2_X1 \myexu/_4986_ ( .A(\myexu/_2344_ ), .B(\myexu/_2280_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1903_ ) );
AND2_X1 \myexu/_4987_ ( .A1(\myexu/_1903_ ), .A2(\myexu/_1838_ ), .ZN(\myexu/_0171_ ) );
NOR2_X1 \myexu/_4988_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2345_ ), .ZN(\myexu/_1904_ ) );
AOI211_X4 \myexu/_4989_ ( .A(\myexu/_2426_ ), .B(\myexu/_1904_ ), .C1(\myexu/_0441_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0172_ ) );
MUX2_X1 \myexu/_4990_ ( .A(\myexu/_2347_ ), .B(\myexu/_2283_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1905_ ) );
AND2_X1 \myexu/_4991_ ( .A1(\myexu/_1905_ ), .A2(\myexu/_2046_ ), .ZN(\myexu/_0173_ ) );
NOR2_X1 \myexu/_4992_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2348_ ), .ZN(\myexu/_1906_ ) );
AOI211_X4 \myexu/_4993_ ( .A(\myexu/_2426_ ), .B(\myexu/_1906_ ), .C1(\myexu/_1544_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0174_ ) );
NOR2_X1 \myexu/_4994_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2531_ ), .ZN(\myexu/_1907_ ) );
AOI211_X4 \myexu/_4995_ ( .A(\myexu/_2426_ ), .B(\myexu/_1907_ ), .C1(\myexu/_2121_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0175_ ) );
NOR2_X1 \myexu/_4996_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2532_ ), .ZN(\myexu/_1908_ ) );
AOI211_X4 \myexu/_4997_ ( .A(\myexu/_2426_ ), .B(\myexu/_1908_ ), .C1(\myexu/_2107_ ), .C2(\myexu/_1895_ ), .ZN(\myexu/_0176_ ) );
NOR2_X1 \myexu/_4998_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2533_ ), .ZN(\myexu/_1909_ ) );
AOI211_X4 \myexu/_4999_ ( .A(\myexu/_2426_ ), .B(\myexu/_1909_ ), .C1(\myexu/_2115_ ), .C2(\myexu/_1987_ ), .ZN(\myexu/_0177_ ) );
NOR2_X1 \myexu/_5000_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2534_ ), .ZN(\myexu/_1910_ ) );
AOI211_X4 \myexu/_5001_ ( .A(\myexu/_2426_ ), .B(\myexu/_1910_ ), .C1(\myexu/_1589_ ), .C2(\myexu/_1987_ ), .ZN(\myexu/_0178_ ) );
NOR2_X1 \myexu/_5002_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_2535_ ), .ZN(\myexu/_1911_ ) );
AOI211_X4 \myexu/_5003_ ( .A(\myexu/_2426_ ), .B(\myexu/_1911_ ), .C1(\myexu/_1939_ ), .C2(\myexu/_1987_ ), .ZN(\myexu/_0179_ ) );
NOR2_X1 \myexu/_5004_ ( .A1(\myexu/_2002_ ), .A2(\myexu/_0292_ ), .ZN(\myexu/_1912_ ) );
AOI211_X4 \myexu/_5005_ ( .A(\myexu/_2426_ ), .B(\myexu/_1912_ ), .C1(\myexu/_2034_ ), .C2(\myexu/_1987_ ), .ZN(\myexu/_0180_ ) );
NOR3_X1 \myexu/_5006_ ( .A1(\myexu/_1970_ ), .A2(\myexu/_2537_ ), .A3(\myexu/_2529_ ), .ZN(\myexu/_1913_ ) );
INV_X1 \myexu/_5007_ ( .A(\myexu/_0293_ ), .ZN(\myexu/_1914_ ) );
AOI211_X4 \myexu/_5008_ ( .A(\myexu/_2426_ ), .B(\myexu/_1913_ ), .C1(\myexu/_1914_ ), .C2(\myexu/_1999_ ), .ZN(\myexu/_0181_ ) );
OAI21_X1 \myexu/_5009_ ( .A(\myexu/_0294_ ), .B1(\myexu/_1970_ ), .B2(\myexu/_2537_ ), .ZN(\myexu/_1915_ ) );
AOI21_X1 \myexu/_5010_ ( .A(\myexu/_2426_ ), .B1(\myexu/_1599_ ), .B2(\myexu/_1915_ ), .ZN(\myexu/_0182_ ) );
MUX2_X1 \myexu/_5011_ ( .A(\myexu/_0287_ ), .B(\myexu/_2356_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1916_ ) );
AND2_X1 \myexu/_5012_ ( .A1(\myexu/_1916_ ), .A2(\myexu/_2046_ ), .ZN(\myexu/_0183_ ) );
MUX2_X1 \myexu/_5013_ ( .A(\myexu/_0288_ ), .B(\myexu/_2357_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1917_ ) );
AND2_X1 \myexu/_5014_ ( .A1(\myexu/_1917_ ), .A2(\myexu/_2046_ ), .ZN(\myexu/_0184_ ) );
MUX2_X1 \myexu/_5015_ ( .A(\myexu/_0289_ ), .B(\myexu/_2358_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1918_ ) );
AND2_X1 \myexu/_5016_ ( .A1(\myexu/_1918_ ), .A2(\myexu/_2046_ ), .ZN(\myexu/_0185_ ) );
MUX2_X1 \myexu/_5017_ ( .A(\myexu/_0290_ ), .B(\myexu/_2359_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1919_ ) );
AND2_X1 \myexu/_5018_ ( .A1(\myexu/_1919_ ), .A2(\myexu/_2046_ ), .ZN(\myexu/_0186_ ) );
MUX2_X1 \myexu/_5019_ ( .A(\myexu/_0291_ ), .B(\myexu/_2360_ ), .S(\myexu/_1891_ ), .Z(\myexu/_1920_ ) );
AND2_X1 \myexu/_5020_ ( .A1(\myexu/_1920_ ), .A2(\myexu/_2046_ ), .ZN(\myexu/_0187_ ) );
NAND2_X1 \myexu/_5021_ ( .A1(\myexu/_1972_ ), .A2(\myexu/_2537_ ), .ZN(\myexu/_1921_ ) );
AOI211_X4 \myexu/_5022_ ( .A(\myexu/_0294_ ), .B(\myexu/_1914_ ), .C1(\myexu/_0000_ ), .C2(\myexu/_0292_ ), .ZN(\myexu/_1922_ ) );
INV_X1 \myexu/_5023_ ( .A(\myexu/_0001_ ), .ZN(\myexu/_1923_ ) );
OAI21_X1 \myexu/_5024_ ( .A(\myexu/_1922_ ), .B1(\myexu/_0292_ ), .B2(\myexu/_1923_ ), .ZN(\myexu/_1924_ ) );
AOI21_X1 \myexu/_5025_ ( .A(\myexu/_1921_ ), .B1(\myexu/_1924_ ), .B2(\myexu/_2361_ ), .ZN(\myexu/_1925_ ) );
OR2_X1 \myexu/_5026_ ( .A1(\myexu/_1925_ ), .A2(\myexu/_1976_ ), .ZN(\myexu/_0188_ ) );
DFF_X1 \myexu/_5027_ ( .D(\myexu/_2712_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(\myexu/_2711_ ) );
DFF_X1 \myexu/_5028_ ( .D(\myexu/_2713_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(\myexu/_2710_ ) );
DFF_X1 \myexu/_5029_ ( .D(\myexu/_2714_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(\myexu/_2709_ ) );
DFF_X1 \myexu/_5030_ ( .D(\myexu/_2715_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(\myexu/_2708_ ) );
DFF_X1 \myexu/_5031_ ( .D(\myexu/_2716_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(\myexu/_2707_ ) );
DFF_X1 \myexu/_5032_ ( .D(\myexu/_2717_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(\myexu/_2706_ ) );
DFF_X1 \myexu/_5033_ ( .D(\myexu/_2718_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(\myexu/_2705_ ) );
DFF_X1 \myexu/_5034_ ( .D(\myexu/_2719_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(\myexu/_2704_ ) );
DFF_X1 \myexu/_5035_ ( .D(\myexu/_2720_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(\myexu/_2703_ ) );
DFF_X1 \myexu/_5036_ ( .D(\myexu/_2721_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(\myexu/_2702_ ) );
DFF_X1 \myexu/_5037_ ( .D(\myexu/_2722_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(\myexu/_2701_ ) );
DFF_X1 \myexu/_5038_ ( .D(\myexu/_2723_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(\myexu/_2700_ ) );
DFF_X1 \myexu/_5039_ ( .D(\myexu/_2724_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(\myexu/_2699_ ) );
DFF_X1 \myexu/_5040_ ( .D(\myexu/_2725_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(\myexu/_2698_ ) );
DFF_X1 \myexu/_5041_ ( .D(\myexu/_2726_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(\myexu/_2697_ ) );
DFF_X1 \myexu/_5042_ ( .D(\myexu/_2727_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(\myexu/_2696_ ) );
DFF_X1 \myexu/_5043_ ( .D(\myexu/_2728_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(\myexu/_2695_ ) );
DFF_X1 \myexu/_5044_ ( .D(\myexu/_2729_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(\myexu/_2694_ ) );
DFF_X1 \myexu/_5045_ ( .D(\myexu/_2730_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(\myexu/_2693_ ) );
DFF_X1 \myexu/_5046_ ( .D(\myexu/_2731_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(\myexu/_2692_ ) );
DFF_X1 \myexu/_5047_ ( .D(\myexu/_2732_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(\myexu/_2691_ ) );
DFF_X1 \myexu/_5048_ ( .D(\myexu/_2733_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(\myexu/_2690_ ) );
DFF_X1 \myexu/_5049_ ( .D(\myexu/_2734_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(\myexu/_2689_ ) );
DFF_X1 \myexu/_5050_ ( .D(\myexu/_2735_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(\myexu/_2688_ ) );
DFF_X1 \myexu/_5051_ ( .D(\myexu/_2736_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(\myexu/_2687_ ) );
DFF_X1 \myexu/_5052_ ( .D(\myexu/_2737_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(\myexu/_2686_ ) );
DFF_X1 \myexu/_5053_ ( .D(\myexu/_2738_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(\myexu/_2685_ ) );
DFF_X1 \myexu/_5054_ ( .D(\myexu/_2739_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(\myexu/_2684_ ) );
DFF_X1 \myexu/_5055_ ( .D(\myexu/_2740_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(\myexu/_2683_ ) );
DFF_X1 \myexu/_5056_ ( .D(\myexu/_2741_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(\myexu/_2682_ ) );
DFF_X1 \myexu/_5057_ ( .D(\myexu/_2742_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(\myexu/_2681_ ) );
DFF_X1 \myexu/_5058_ ( .D(\myexu/_2743_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(\myexu/_2680_ ) );
DFF_X1 \myexu/_5059_ ( .D(\myexu/_2744_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(\myexu/_2679_ ) );
DFF_X1 \myexu/_5060_ ( .D(\myexu/_2745_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(\myexu/_2678_ ) );
DFF_X1 \myexu/_5061_ ( .D(\myexu/_2746_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(\myexu/_2677_ ) );
DFF_X1 \myexu/_5062_ ( .D(\myexu/_2747_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(\myexu/_2676_ ) );
DFF_X1 \myexu/_5063_ ( .D(\myexu/_2748_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(\myexu/_2675_ ) );
DFF_X1 \myexu/_5064_ ( .D(\myexu/_2749_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(\myexu/_2674_ ) );
DFF_X1 \myexu/_5065_ ( .D(\myexu/_2750_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(\myexu/_2673_ ) );
DFF_X1 \myexu/_5066_ ( .D(\myexu/_2751_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(\myexu/_2672_ ) );
DFF_X1 \myexu/_5067_ ( .D(\myexu/_2752_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(\myexu/_2671_ ) );
DFF_X1 \myexu/_5068_ ( .D(\myexu/_2753_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(\myexu/_2670_ ) );
DFF_X1 \myexu/_5069_ ( .D(\myexu/_2754_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(\myexu/_2669_ ) );
DFF_X1 \myexu/_5070_ ( .D(\myexu/_2755_ ), .CK(clock ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(\myexu/_2668_ ) );
DFF_X1 \myexu/_5071_ ( .D(\myexu/_2756_ ), .CK(clock ), .Q(\pc_jump [0] ), .QN(\myexu/_2667_ ) );
DFF_X1 \myexu/_5072_ ( .D(\myexu/_2757_ ), .CK(clock ), .Q(\pc_jump [1] ), .QN(\myexu/_2666_ ) );
DFF_X1 \myexu/_5073_ ( .D(\myexu/_2758_ ), .CK(clock ), .Q(\pc_jump [2] ), .QN(\myexu/_2665_ ) );
DFF_X1 \myexu/_5074_ ( .D(\myexu/_2759_ ), .CK(clock ), .Q(\pc_jump [3] ), .QN(\myexu/_2664_ ) );
DFF_X1 \myexu/_5075_ ( .D(\myexu/_2760_ ), .CK(clock ), .Q(\pc_jump [4] ), .QN(\myexu/_2663_ ) );
DFF_X1 \myexu/_5076_ ( .D(\myexu/_2761_ ), .CK(clock ), .Q(\pc_jump [5] ), .QN(\myexu/_2662_ ) );
DFF_X1 \myexu/_5077_ ( .D(\myexu/_2762_ ), .CK(clock ), .Q(\pc_jump [6] ), .QN(\myexu/_2661_ ) );
DFF_X1 \myexu/_5078_ ( .D(\myexu/_2763_ ), .CK(clock ), .Q(\pc_jump [7] ), .QN(\myexu/_2660_ ) );
DFF_X1 \myexu/_5079_ ( .D(\myexu/_2764_ ), .CK(clock ), .Q(\pc_jump [8] ), .QN(\myexu/_2659_ ) );
DFF_X1 \myexu/_5080_ ( .D(\myexu/_2765_ ), .CK(clock ), .Q(\pc_jump [9] ), .QN(\myexu/_2658_ ) );
DFF_X1 \myexu/_5081_ ( .D(\myexu/_2766_ ), .CK(clock ), .Q(\pc_jump [10] ), .QN(\myexu/_2657_ ) );
DFF_X1 \myexu/_5082_ ( .D(\myexu/_2767_ ), .CK(clock ), .Q(\pc_jump [11] ), .QN(\myexu/_2656_ ) );
DFF_X1 \myexu/_5083_ ( .D(\myexu/_2768_ ), .CK(clock ), .Q(\pc_jump [12] ), .QN(\myexu/_2655_ ) );
DFF_X1 \myexu/_5084_ ( .D(\myexu/_2769_ ), .CK(clock ), .Q(\pc_jump [13] ), .QN(\myexu/_2654_ ) );
DFF_X1 \myexu/_5085_ ( .D(\myexu/_2770_ ), .CK(clock ), .Q(\pc_jump [14] ), .QN(\myexu/_2653_ ) );
DFF_X1 \myexu/_5086_ ( .D(\myexu/_2771_ ), .CK(clock ), .Q(\pc_jump [15] ), .QN(\myexu/_2652_ ) );
DFF_X1 \myexu/_5087_ ( .D(\myexu/_2772_ ), .CK(clock ), .Q(\pc_jump [16] ), .QN(\myexu/_2651_ ) );
DFF_X1 \myexu/_5088_ ( .D(\myexu/_2773_ ), .CK(clock ), .Q(\pc_jump [17] ), .QN(\myexu/_2650_ ) );
DFF_X1 \myexu/_5089_ ( .D(\myexu/_2774_ ), .CK(clock ), .Q(\pc_jump [18] ), .QN(\myexu/_2649_ ) );
DFF_X1 \myexu/_5090_ ( .D(\myexu/_2775_ ), .CK(clock ), .Q(\pc_jump [19] ), .QN(\myexu/_2648_ ) );
DFF_X1 \myexu/_5091_ ( .D(\myexu/_2776_ ), .CK(clock ), .Q(\pc_jump [20] ), .QN(\myexu/_2647_ ) );
DFF_X1 \myexu/_5092_ ( .D(\myexu/_2777_ ), .CK(clock ), .Q(\pc_jump [21] ), .QN(\myexu/_2646_ ) );
DFF_X1 \myexu/_5093_ ( .D(\myexu/_2778_ ), .CK(clock ), .Q(\pc_jump [22] ), .QN(\myexu/_2645_ ) );
DFF_X1 \myexu/_5094_ ( .D(\myexu/_2779_ ), .CK(clock ), .Q(\pc_jump [23] ), .QN(\myexu/_2644_ ) );
DFF_X1 \myexu/_5095_ ( .D(\myexu/_2780_ ), .CK(clock ), .Q(\pc_jump [24] ), .QN(\myexu/_2643_ ) );
DFF_X1 \myexu/_5096_ ( .D(\myexu/_2781_ ), .CK(clock ), .Q(\pc_jump [25] ), .QN(\myexu/_2642_ ) );
DFF_X1 \myexu/_5097_ ( .D(\myexu/_2782_ ), .CK(clock ), .Q(\pc_jump [26] ), .QN(\myexu/_2641_ ) );
DFF_X1 \myexu/_5098_ ( .D(\myexu/_2783_ ), .CK(clock ), .Q(\pc_jump [27] ), .QN(\myexu/_2640_ ) );
DFF_X1 \myexu/_5099_ ( .D(\myexu/_2784_ ), .CK(clock ), .Q(\pc_jump [28] ), .QN(\myexu/_2639_ ) );
DFF_X1 \myexu/_5100_ ( .D(\myexu/_2785_ ), .CK(clock ), .Q(\pc_jump [29] ), .QN(\myexu/_2638_ ) );
DFF_X1 \myexu/_5101_ ( .D(\myexu/_2786_ ), .CK(clock ), .Q(\pc_jump [30] ), .QN(\myexu/_2637_ ) );
DFF_X1 \myexu/_5102_ ( .D(\myexu/_2787_ ), .CK(clock ), .Q(\pc_jump [31] ), .QN(\myexu/_2636_ ) );
DFF_X1 \myexu/_5103_ ( .D(\myexu/_2788_ ), .CK(clock ), .Q(check_quest ), .QN(\myexu/_2635_ ) );
DFF_X1 \myexu/_5104_ ( .D(\myexu/_2789_ ), .CK(clock ), .Q(\EX_LS_pc [0] ), .QN(\myexu/_2634_ ) );
DFF_X1 \myexu/_5105_ ( .D(\myexu/_2790_ ), .CK(clock ), .Q(\EX_LS_pc [1] ), .QN(\myexu/_2633_ ) );
DFF_X1 \myexu/_5106_ ( .D(\myexu/_2791_ ), .CK(clock ), .Q(\EX_LS_pc [2] ), .QN(\myexu/_2632_ ) );
DFF_X1 \myexu/_5107_ ( .D(\myexu/_2792_ ), .CK(clock ), .Q(\EX_LS_pc [3] ), .QN(\myexu/_2631_ ) );
DFF_X1 \myexu/_5108_ ( .D(\myexu/_2793_ ), .CK(clock ), .Q(\EX_LS_pc [4] ), .QN(\myexu/_2630_ ) );
DFF_X1 \myexu/_5109_ ( .D(\myexu/_2794_ ), .CK(clock ), .Q(\EX_LS_pc [5] ), .QN(\myexu/_2629_ ) );
DFF_X1 \myexu/_5110_ ( .D(\myexu/_2795_ ), .CK(clock ), .Q(\EX_LS_pc [6] ), .QN(\myexu/_2628_ ) );
DFF_X1 \myexu/_5111_ ( .D(\myexu/_2796_ ), .CK(clock ), .Q(\EX_LS_pc [7] ), .QN(\myexu/_2627_ ) );
DFF_X1 \myexu/_5112_ ( .D(\myexu/_2797_ ), .CK(clock ), .Q(\EX_LS_pc [8] ), .QN(\myexu/_2626_ ) );
DFF_X1 \myexu/_5113_ ( .D(\myexu/_2798_ ), .CK(clock ), .Q(\EX_LS_pc [9] ), .QN(\myexu/_2625_ ) );
DFF_X1 \myexu/_5114_ ( .D(\myexu/_2799_ ), .CK(clock ), .Q(\EX_LS_pc [10] ), .QN(\myexu/_2624_ ) );
DFF_X1 \myexu/_5115_ ( .D(\myexu/_2800_ ), .CK(clock ), .Q(\EX_LS_pc [11] ), .QN(\myexu/_2623_ ) );
DFF_X1 \myexu/_5116_ ( .D(\myexu/_2801_ ), .CK(clock ), .Q(\EX_LS_pc [12] ), .QN(\myexu/_2622_ ) );
DFF_X1 \myexu/_5117_ ( .D(\myexu/_2802_ ), .CK(clock ), .Q(\EX_LS_pc [13] ), .QN(\myexu/_2621_ ) );
DFF_X1 \myexu/_5118_ ( .D(\myexu/_2803_ ), .CK(clock ), .Q(\EX_LS_pc [14] ), .QN(\myexu/_2620_ ) );
DFF_X1 \myexu/_5119_ ( .D(\myexu/_2804_ ), .CK(clock ), .Q(\EX_LS_pc [15] ), .QN(\myexu/_2619_ ) );
DFF_X1 \myexu/_5120_ ( .D(\myexu/_2805_ ), .CK(clock ), .Q(\EX_LS_pc [16] ), .QN(\myexu/_2618_ ) );
DFF_X1 \myexu/_5121_ ( .D(\myexu/_2806_ ), .CK(clock ), .Q(\EX_LS_pc [17] ), .QN(\myexu/_2617_ ) );
DFF_X1 \myexu/_5122_ ( .D(\myexu/_2807_ ), .CK(clock ), .Q(\EX_LS_pc [18] ), .QN(\myexu/_2616_ ) );
DFF_X1 \myexu/_5123_ ( .D(\myexu/_2808_ ), .CK(clock ), .Q(\EX_LS_pc [19] ), .QN(\myexu/_2615_ ) );
DFF_X1 \myexu/_5124_ ( .D(\myexu/_2809_ ), .CK(clock ), .Q(\EX_LS_pc [20] ), .QN(\myexu/_2614_ ) );
DFF_X1 \myexu/_5125_ ( .D(\myexu/_2810_ ), .CK(clock ), .Q(\EX_LS_pc [21] ), .QN(\myexu/_2613_ ) );
DFF_X1 \myexu/_5126_ ( .D(\myexu/_2811_ ), .CK(clock ), .Q(\EX_LS_pc [22] ), .QN(\myexu/_2612_ ) );
DFF_X1 \myexu/_5127_ ( .D(\myexu/_2812_ ), .CK(clock ), .Q(\EX_LS_pc [23] ), .QN(\myexu/_2611_ ) );
DFF_X1 \myexu/_5128_ ( .D(\myexu/_2813_ ), .CK(clock ), .Q(\EX_LS_pc [24] ), .QN(\myexu/_2610_ ) );
DFF_X1 \myexu/_5129_ ( .D(\myexu/_2814_ ), .CK(clock ), .Q(\EX_LS_pc [25] ), .QN(\myexu/_2609_ ) );
DFF_X1 \myexu/_5130_ ( .D(\myexu/_2815_ ), .CK(clock ), .Q(\EX_LS_pc [26] ), .QN(\myexu/_2608_ ) );
DFF_X1 \myexu/_5131_ ( .D(\myexu/_2816_ ), .CK(clock ), .Q(\EX_LS_pc [27] ), .QN(\myexu/_2607_ ) );
DFF_X1 \myexu/_5132_ ( .D(\myexu/_2817_ ), .CK(clock ), .Q(\EX_LS_pc [28] ), .QN(\myexu/_2606_ ) );
DFF_X1 \myexu/_5133_ ( .D(\myexu/_2818_ ), .CK(clock ), .Q(\EX_LS_pc [29] ), .QN(\myexu/_2605_ ) );
DFF_X1 \myexu/_5134_ ( .D(\myexu/_2819_ ), .CK(clock ), .Q(\EX_LS_pc [30] ), .QN(\myexu/_2604_ ) );
DFF_X1 \myexu/_5135_ ( .D(\myexu/_2820_ ), .CK(clock ), .Q(\EX_LS_pc [31] ), .QN(\myexu/_2603_ ) );
DFF_X1 \myexu/_5136_ ( .D(\myexu/_2821_ ), .CK(clock ), .Q(\EX_LS_typ [0] ), .QN(\myexu/_2602_ ) );
DFF_X1 \myexu/_5137_ ( .D(\myexu/_2822_ ), .CK(clock ), .Q(\EX_LS_typ [1] ), .QN(\myexu/_2601_ ) );
DFF_X1 \myexu/_5138_ ( .D(\myexu/_2823_ ), .CK(clock ), .Q(\EX_LS_typ [2] ), .QN(\myexu/_2600_ ) );
DFF_X1 \myexu/_5139_ ( .D(\myexu/_2824_ ), .CK(clock ), .Q(\EX_LS_typ [3] ), .QN(\myexu/_2599_ ) );
DFF_X1 \myexu/_5140_ ( .D(\myexu/_2825_ ), .CK(clock ), .Q(\EX_LS_typ [4] ), .QN(\myexu/_2598_ ) );
DFF_X1 \myexu/_5141_ ( .D(\myexu/_2826_ ), .CK(clock ), .Q(\EX_LS_flag [0] ), .QN(\myexu/_2597_ ) );
DFF_X1 \myexu/_5142_ ( .D(\myexu/_2827_ ), .CK(clock ), .Q(\EX_LS_flag [1] ), .QN(\myexu/_2596_ ) );
DFF_X1 \myexu/_5143_ ( .D(\myexu/_2828_ ), .CK(clock ), .Q(\EX_LS_flag [2] ), .QN(\myexu/_2595_ ) );
DFF_X1 \myexu/_5144_ ( .D(\myexu/_2829_ ), .CK(clock ), .Q(\EX_LS_dest_reg [0] ), .QN(\myexu/_2594_ ) );
DFF_X1 \myexu/_5145_ ( .D(\myexu/_2830_ ), .CK(clock ), .Q(\EX_LS_dest_reg [1] ), .QN(\myexu/_2593_ ) );
DFF_X1 \myexu/_5146_ ( .D(\myexu/_2831_ ), .CK(clock ), .Q(\EX_LS_dest_reg [2] ), .QN(\myexu/_2592_ ) );
DFF_X1 \myexu/_5147_ ( .D(\myexu/_2832_ ), .CK(clock ), .Q(\EX_LS_dest_reg [3] ), .QN(\myexu/_2591_ ) );
DFF_X1 \myexu/_5148_ ( .D(\myexu/_2833_ ), .CK(clock ), .Q(\EX_LS_dest_reg [4] ), .QN(\myexu/_2590_ ) );
DFF_X1 \myexu/_5149_ ( .D(\myexu/_2834_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(EXU_ready_IDU ) );
DFF_X1 \myexu/_5150_ ( .D(\myexu/_2835_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(\myexu/_2589_ ) );
DFF_X1 \myexu/_5151_ ( .D(\myexu/_2836_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(\myexu/_2588_ ) );
DFF_X1 \myexu/_5152_ ( .D(\myexu/_2837_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(\myexu/_2587_ ) );
DFF_X1 \myexu/_5153_ ( .D(\myexu/_2838_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(\myexu/_2586_ ) );
DFF_X1 \myexu/_5154_ ( .D(\myexu/_2839_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(\myexu/_2585_ ) );
DFF_X1 \myexu/_5155_ ( .D(\myexu/_2840_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(\myexu/_2584_ ) );
DFF_X1 \myexu/_5156_ ( .D(\myexu/_2841_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(\myexu/_2583_ ) );
DFF_X1 \myexu/_5157_ ( .D(\myexu/_2842_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(\myexu/_2582_ ) );
DFF_X1 \myexu/_5158_ ( .D(\myexu/_2843_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(\myexu/_2581_ ) );
DFF_X1 \myexu/_5159_ ( .D(\myexu/_2844_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(\myexu/_2580_ ) );
DFF_X1 \myexu/_5160_ ( .D(\myexu/_2845_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(\myexu/_2579_ ) );
DFF_X1 \myexu/_5161_ ( .D(\myexu/_2846_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(\myexu/_2578_ ) );
DFF_X1 \myexu/_5162_ ( .D(\myexu/_2847_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(\myexu/_2577_ ) );
DFF_X1 \myexu/_5163_ ( .D(\myexu/_2848_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(\myexu/_2576_ ) );
DFF_X1 \myexu/_5164_ ( .D(\myexu/_2849_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(\myexu/_2575_ ) );
DFF_X1 \myexu/_5165_ ( .D(\myexu/_2850_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(\myexu/_2574_ ) );
DFF_X1 \myexu/_5166_ ( .D(\myexu/_2851_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(\myexu/_2573_ ) );
DFF_X1 \myexu/_5167_ ( .D(\myexu/_2852_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(\myexu/_2572_ ) );
DFF_X1 \myexu/_5168_ ( .D(\myexu/_2853_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(\myexu/_2571_ ) );
DFF_X1 \myexu/_5169_ ( .D(\myexu/_2854_ ), .CK(clock ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(\myexu/_2570_ ) );
DFF_X1 \myexu/_5170_ ( .D(\myexu/_2855_ ), .CK(clock ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu/_2569_ ) );
DFF_X1 \myexu/_5171_ ( .D(\myexu/_2856_ ), .CK(clock ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu/_2568_ ) );
DFF_X1 \myexu/_5172_ ( .D(\myexu/_2857_ ), .CK(clock ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu/_2567_ ) );
DFF_X1 \myexu/_5173_ ( .D(\myexu/_2858_ ), .CK(clock ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu/_2566_ ) );
DFF_X1 \myexu/_5174_ ( .D(\myexu/_2859_ ), .CK(clock ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu/_2565_ ) );
DFF_X1 \myexu/_5175_ ( .D(\myexu/_2860_ ), .CK(clock ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu/_2564_ ) );
DFF_X1 \myexu/_5176_ ( .D(\myexu/_2861_ ), .CK(clock ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu/_2563_ ) );
DFF_X1 \myexu/_5177_ ( .D(\myexu/_2862_ ), .CK(clock ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu/_2562_ ) );
DFF_X1 \myexu/_5178_ ( .D(\myexu/_2863_ ), .CK(clock ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu/_2561_ ) );
DFF_X1 \myexu/_5179_ ( .D(\myexu/_2864_ ), .CK(clock ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu/_2560_ ) );
DFF_X1 \myexu/_5180_ ( .D(\myexu/_2865_ ), .CK(clock ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu/_2559_ ) );
DFF_X1 \myexu/_5181_ ( .D(\myexu/_2866_ ), .CK(clock ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu/_2558_ ) );
DFF_X1 \myexu/_5182_ ( .D(\myexu/_2867_ ), .CK(clock ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu/_2557_ ) );
DFF_X1 \myexu/_5183_ ( .D(\myexu/_2868_ ), .CK(clock ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu/_2556_ ) );
DFF_X1 \myexu/_5184_ ( .D(\myexu/_2869_ ), .CK(clock ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu/_2555_ ) );
DFF_X1 \myexu/_5185_ ( .D(\myexu/_2870_ ), .CK(clock ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu/_2554_ ) );
DFF_X1 \myexu/_5186_ ( .D(\myexu/_2871_ ), .CK(clock ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu/_2553_ ) );
DFF_X1 \myexu/_5187_ ( .D(\myexu/_2872_ ), .CK(clock ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu/_2552_ ) );
DFF_X1 \myexu/_5188_ ( .D(\myexu/_2873_ ), .CK(clock ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu/_2551_ ) );
DFF_X1 \myexu/_5189_ ( .D(\myexu/_2874_ ), .CK(clock ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu/_2550_ ) );
DFF_X1 \myexu/_5190_ ( .D(\myexu/_2875_ ), .CK(clock ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu/_2549_ ) );
DFF_X1 \myexu/_5191_ ( .D(\myexu/_2876_ ), .CK(clock ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu/_2548_ ) );
DFF_X1 \myexu/_5192_ ( .D(\myexu/_2877_ ), .CK(clock ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu/_2547_ ) );
DFF_X1 \myexu/_5193_ ( .D(\myexu/_2878_ ), .CK(clock ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu/_2546_ ) );
DFF_X1 \myexu/_5194_ ( .D(\myexu/_2879_ ), .CK(clock ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu/_2545_ ) );
DFF_X1 \myexu/_5195_ ( .D(\myexu/_2880_ ), .CK(clock ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu/_2544_ ) );
DFF_X1 \myexu/_5196_ ( .D(\myexu/_2881_ ), .CK(clock ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu/_2543_ ) );
DFF_X1 \myexu/_5197_ ( .D(\myexu/_2882_ ), .CK(clock ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu/_2542_ ) );
DFF_X1 \myexu/_5198_ ( .D(\myexu/_2883_ ), .CK(clock ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu/_2541_ ) );
DFF_X1 \myexu/_5199_ ( .D(\myexu/_2884_ ), .CK(clock ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu/_2540_ ) );
DFF_X1 \myexu/_5200_ ( .D(\myexu/_2885_ ), .CK(clock ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu/_2539_ ) );
DFF_X1 \myexu/_5201_ ( .D(\myexu/_2886_ ), .CK(clock ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu/_2538_ ) );
BUF_X1 \myexu/_5202_ ( .A(\EX_LS_flag [0] ), .Z(\EX_LS_typ [5] ) );
BUF_X1 \myexu/_5203_ ( .A(\EX_LS_flag [1] ), .Z(\EX_LS_typ [6] ) );
BUF_X1 \myexu/_5204_ ( .A(\EX_LS_flag [2] ), .Z(\EX_LS_typ [7] ) );
BUF_X1 \myexu/_5205_ ( .A(\src2 [31] ), .Z(\myexu/_2483_ ) );
BUF_X1 \myexu/_5206_ ( .A(\ID_EX_imm [31] ), .Z(\myexu/_0319_ ) );
BUF_X1 \myexu/_5207_ ( .A(\ID_EX_typ [4] ), .Z(\myexu/_2527_ ) );
BUF_X1 \myexu/_5208_ ( .A(\myexu/_0026_ ), .Z(\myexu/alu_op [31] ) );
BUF_X1 \myexu/_5209_ ( .A(\src1 [12] ), .Z(\myexu/_2430_ ) );
BUF_X1 \myexu/_5210_ ( .A(\ID_EX_imm [12] ), .Z(\myexu/_0298_ ) );
BUF_X1 \myexu/_5211_ ( .A(\src1 [11] ), .Z(\myexu/_2429_ ) );
BUF_X1 \myexu/_5212_ ( .A(\ID_EX_imm [11] ), .Z(\myexu/_0297_ ) );
BUF_X1 \myexu/_5213_ ( .A(\src1 [10] ), .Z(\myexu/_2428_ ) );
BUF_X1 \myexu/_5214_ ( .A(\ID_EX_imm [10] ), .Z(\myexu/_0296_ ) );
BUF_X1 \myexu/_5215_ ( .A(\src1 [9] ), .Z(\myexu/_2458_ ) );
BUF_X1 \myexu/_5216_ ( .A(\ID_EX_imm [9] ), .Z(\myexu/_0326_ ) );
BUF_X1 \myexu/_5217_ ( .A(\src1 [8] ), .Z(\myexu/_2457_ ) );
BUF_X1 \myexu/_5218_ ( .A(\ID_EX_imm [8] ), .Z(\myexu/_0325_ ) );
BUF_X1 \myexu/_5219_ ( .A(\src1 [7] ), .Z(\myexu/_2456_ ) );
BUF_X1 \myexu/_5220_ ( .A(\ID_EX_imm [7] ), .Z(\myexu/_0324_ ) );
BUF_X1 \myexu/_5221_ ( .A(\src1 [6] ), .Z(\myexu/_2455_ ) );
BUF_X1 \myexu/_5222_ ( .A(\ID_EX_imm [6] ), .Z(\myexu/_0323_ ) );
BUF_X1 \myexu/_5223_ ( .A(\src1 [5] ), .Z(\myexu/_2454_ ) );
BUF_X1 \myexu/_5224_ ( .A(\ID_EX_imm [5] ), .Z(\myexu/_0322_ ) );
BUF_X1 \myexu/_5225_ ( .A(\src1 [4] ), .Z(\myexu/_2453_ ) );
BUF_X1 \myexu/_5226_ ( .A(\ID_EX_imm [4] ), .Z(\myexu/_0321_ ) );
BUF_X1 \myexu/_5227_ ( .A(\src1 [3] ), .Z(\myexu/_2452_ ) );
BUF_X1 \myexu/_5228_ ( .A(\ID_EX_imm [3] ), .Z(\myexu/_0320_ ) );
BUF_X1 \myexu/_5229_ ( .A(\src1 [2] ), .Z(\myexu/_2449_ ) );
BUF_X1 \myexu/_5230_ ( .A(\ID_EX_imm [2] ), .Z(\myexu/_0317_ ) );
BUF_X1 \myexu/_5231_ ( .A(\src1 [1] ), .Z(\myexu/_2438_ ) );
BUF_X1 \myexu/_5232_ ( .A(\ID_EX_imm [1] ), .Z(\myexu/_0306_ ) );
BUF_X1 \myexu/_5233_ ( .A(\src1 [0] ), .Z(\myexu/_2427_ ) );
BUF_X1 \myexu/_5234_ ( .A(\ID_EX_imm [0] ), .Z(\myexu/_0295_ ) );
BUF_X1 \myexu/_5235_ ( .A(\src1 [13] ), .Z(\myexu/_2431_ ) );
BUF_X1 \myexu/_5236_ ( .A(\ID_EX_imm [13] ), .Z(\myexu/_0299_ ) );
BUF_X1 \myexu/_5237_ ( .A(\src1 [14] ), .Z(\myexu/_2432_ ) );
BUF_X1 \myexu/_5238_ ( .A(\ID_EX_imm [14] ), .Z(\myexu/_0300_ ) );
BUF_X1 \myexu/_5239_ ( .A(\src1 [15] ), .Z(\myexu/_2433_ ) );
BUF_X1 \myexu/_5240_ ( .A(\ID_EX_imm [15] ), .Z(\myexu/_0301_ ) );
BUF_X1 \myexu/_5241_ ( .A(\src1 [16] ), .Z(\myexu/_2434_ ) );
BUF_X1 \myexu/_5242_ ( .A(\ID_EX_imm [16] ), .Z(\myexu/_0302_ ) );
BUF_X1 \myexu/_5243_ ( .A(\src1 [17] ), .Z(\myexu/_2435_ ) );
BUF_X1 \myexu/_5244_ ( .A(\ID_EX_imm [17] ), .Z(\myexu/_0303_ ) );
BUF_X1 \myexu/_5245_ ( .A(\src1 [18] ), .Z(\myexu/_2436_ ) );
BUF_X1 \myexu/_5246_ ( .A(\ID_EX_imm [18] ), .Z(\myexu/_0304_ ) );
BUF_X1 \myexu/_5247_ ( .A(\src1 [19] ), .Z(\myexu/_2437_ ) );
BUF_X1 \myexu/_5248_ ( .A(\ID_EX_imm [19] ), .Z(\myexu/_0305_ ) );
BUF_X1 \myexu/_5249_ ( .A(\src1 [20] ), .Z(\myexu/_2439_ ) );
BUF_X1 \myexu/_5250_ ( .A(\ID_EX_imm [20] ), .Z(\myexu/_0307_ ) );
BUF_X1 \myexu/_5251_ ( .A(\src1 [21] ), .Z(\myexu/_2440_ ) );
BUF_X1 \myexu/_5252_ ( .A(\ID_EX_imm [21] ), .Z(\myexu/_0308_ ) );
BUF_X1 \myexu/_5253_ ( .A(\src1 [22] ), .Z(\myexu/_2441_ ) );
BUF_X1 \myexu/_5254_ ( .A(\ID_EX_imm [22] ), .Z(\myexu/_0309_ ) );
BUF_X1 \myexu/_5255_ ( .A(\src1 [23] ), .Z(\myexu/_2442_ ) );
BUF_X1 \myexu/_5256_ ( .A(\ID_EX_imm [23] ), .Z(\myexu/_0310_ ) );
BUF_X1 \myexu/_5257_ ( .A(\src1 [24] ), .Z(\myexu/_2443_ ) );
BUF_X1 \myexu/_5258_ ( .A(\ID_EX_imm [24] ), .Z(\myexu/_0311_ ) );
BUF_X1 \myexu/_5259_ ( .A(\src1 [25] ), .Z(\myexu/_2444_ ) );
BUF_X1 \myexu/_5260_ ( .A(\ID_EX_imm [25] ), .Z(\myexu/_0312_ ) );
BUF_X1 \myexu/_5261_ ( .A(\src1 [26] ), .Z(\myexu/_2445_ ) );
BUF_X1 \myexu/_5262_ ( .A(\ID_EX_imm [26] ), .Z(\myexu/_0313_ ) );
BUF_X1 \myexu/_5263_ ( .A(\src1 [27] ), .Z(\myexu/_2446_ ) );
BUF_X1 \myexu/_5264_ ( .A(\ID_EX_imm [27] ), .Z(\myexu/_0314_ ) );
BUF_X1 \myexu/_5265_ ( .A(\src1 [28] ), .Z(\myexu/_2447_ ) );
BUF_X1 \myexu/_5266_ ( .A(\ID_EX_imm [28] ), .Z(\myexu/_0315_ ) );
BUF_X1 \myexu/_5267_ ( .A(\src1 [29] ), .Z(\myexu/_2448_ ) );
BUF_X1 \myexu/_5268_ ( .A(\ID_EX_imm [29] ), .Z(\myexu/_0316_ ) );
BUF_X1 \myexu/_5269_ ( .A(\src1 [30] ), .Z(\myexu/_2450_ ) );
BUF_X1 \myexu/_5270_ ( .A(\ID_EX_imm [30] ), .Z(\myexu/_0318_ ) );
BUF_X1 \myexu/_5271_ ( .A(\src1 [31] ), .Z(\myexu/_2451_ ) );
BUF_X1 \myexu/_5272_ ( .A(IDU_valid_EXU ), .Z(\myexu/_2536_ ) );
BUF_X1 \myexu/_5273_ ( .A(EXU_valid_LSU ), .Z(\myexu/_2537_ ) );
BUF_X1 \myexu/_5274_ ( .A(reset ), .Z(\myexu/_2426_ ) );
BUF_X1 \myexu/_5275_ ( .A(\ID_EX_typ [5] ), .Z(\myexu/_2528_ ) );
BUF_X1 \myexu/_5276_ ( .A(\ID_EX_typ [6] ), .Z(\myexu/_2529_ ) );
BUF_X1 \myexu/_5277_ ( .A(\ID_EX_typ [7] ), .Z(\myexu/_2530_ ) );
BUF_X1 \myexu/_5278_ ( .A(\src2 [0] ), .Z(\myexu/_2459_ ) );
BUF_X1 \myexu/_5279_ ( .A(\myexu/_0002_ ), .Z(\myexu/alu_op [0] ) );
BUF_X1 \myexu/_5280_ ( .A(\src2 [1] ), .Z(\myexu/_2470_ ) );
BUF_X1 \myexu/_5281_ ( .A(\myexu/_0013_ ), .Z(\myexu/alu_op [1] ) );
BUF_X1 \myexu/_5282_ ( .A(\src2 [2] ), .Z(\myexu/_2481_ ) );
BUF_X1 \myexu/_5283_ ( .A(\myexu/_0024_ ), .Z(\myexu/alu_op [2] ) );
BUF_X1 \myexu/_5284_ ( .A(\src2 [3] ), .Z(\myexu/_2484_ ) );
BUF_X1 \myexu/_5285_ ( .A(\myexu/_0027_ ), .Z(\myexu/alu_op [3] ) );
BUF_X1 \myexu/_5286_ ( .A(\src2 [4] ), .Z(\myexu/_2485_ ) );
BUF_X1 \myexu/_5287_ ( .A(\myexu/_0028_ ), .Z(\myexu/alu_op [4] ) );
BUF_X1 \myexu/_5288_ ( .A(\src2 [5] ), .Z(\myexu/_2486_ ) );
BUF_X1 \myexu/_5289_ ( .A(\myexu/_0029_ ), .Z(\myexu/alu_op [5] ) );
BUF_X1 \myexu/_5290_ ( .A(\src2 [6] ), .Z(\myexu/_2487_ ) );
BUF_X1 \myexu/_5291_ ( .A(\myexu/_0030_ ), .Z(\myexu/alu_op [6] ) );
BUF_X1 \myexu/_5292_ ( .A(\src2 [7] ), .Z(\myexu/_2488_ ) );
BUF_X1 \myexu/_5293_ ( .A(\myexu/_0031_ ), .Z(\myexu/alu_op [7] ) );
BUF_X1 \myexu/_5294_ ( .A(\src2 [8] ), .Z(\myexu/_2489_ ) );
BUF_X1 \myexu/_5295_ ( .A(\myexu/_0032_ ), .Z(\myexu/alu_op [8] ) );
BUF_X1 \myexu/_5296_ ( .A(\src2 [9] ), .Z(\myexu/_2490_ ) );
BUF_X1 \myexu/_5297_ ( .A(\myexu/_0033_ ), .Z(\myexu/alu_op [9] ) );
BUF_X1 \myexu/_5298_ ( .A(\src2 [10] ), .Z(\myexu/_2460_ ) );
BUF_X1 \myexu/_5299_ ( .A(\myexu/_0003_ ), .Z(\myexu/alu_op [10] ) );
BUF_X1 \myexu/_5300_ ( .A(\src2 [11] ), .Z(\myexu/_2461_ ) );
BUF_X1 \myexu/_5301_ ( .A(\myexu/_0004_ ), .Z(\myexu/alu_op [11] ) );
BUF_X1 \myexu/_5302_ ( .A(\src2 [12] ), .Z(\myexu/_2462_ ) );
BUF_X1 \myexu/_5303_ ( .A(\myexu/_0005_ ), .Z(\myexu/alu_op [12] ) );
BUF_X1 \myexu/_5304_ ( .A(\src2 [13] ), .Z(\myexu/_2463_ ) );
BUF_X1 \myexu/_5305_ ( .A(\myexu/_0006_ ), .Z(\myexu/alu_op [13] ) );
BUF_X1 \myexu/_5306_ ( .A(\src2 [14] ), .Z(\myexu/_2464_ ) );
BUF_X1 \myexu/_5307_ ( .A(\myexu/_0007_ ), .Z(\myexu/alu_op [14] ) );
BUF_X1 \myexu/_5308_ ( .A(\src2 [15] ), .Z(\myexu/_2465_ ) );
BUF_X1 \myexu/_5309_ ( .A(\myexu/_0008_ ), .Z(\myexu/alu_op [15] ) );
BUF_X1 \myexu/_5310_ ( .A(\src2 [16] ), .Z(\myexu/_2466_ ) );
BUF_X1 \myexu/_5311_ ( .A(\myexu/_0009_ ), .Z(\myexu/alu_op [16] ) );
BUF_X1 \myexu/_5312_ ( .A(\src2 [17] ), .Z(\myexu/_2467_ ) );
BUF_X1 \myexu/_5313_ ( .A(\myexu/_0010_ ), .Z(\myexu/alu_op [17] ) );
BUF_X1 \myexu/_5314_ ( .A(\src2 [18] ), .Z(\myexu/_2468_ ) );
BUF_X1 \myexu/_5315_ ( .A(\myexu/_0011_ ), .Z(\myexu/alu_op [18] ) );
BUF_X1 \myexu/_5316_ ( .A(\src2 [19] ), .Z(\myexu/_2469_ ) );
BUF_X1 \myexu/_5317_ ( .A(\myexu/_0012_ ), .Z(\myexu/alu_op [19] ) );
BUF_X1 \myexu/_5318_ ( .A(\src2 [20] ), .Z(\myexu/_2471_ ) );
BUF_X1 \myexu/_5319_ ( .A(\myexu/_0014_ ), .Z(\myexu/alu_op [20] ) );
BUF_X1 \myexu/_5320_ ( .A(\src2 [21] ), .Z(\myexu/_2472_ ) );
BUF_X1 \myexu/_5321_ ( .A(\myexu/_0015_ ), .Z(\myexu/alu_op [21] ) );
BUF_X1 \myexu/_5322_ ( .A(\src2 [22] ), .Z(\myexu/_2473_ ) );
BUF_X1 \myexu/_5323_ ( .A(\myexu/_0016_ ), .Z(\myexu/alu_op [22] ) );
BUF_X1 \myexu/_5324_ ( .A(\src2 [23] ), .Z(\myexu/_2474_ ) );
BUF_X1 \myexu/_5325_ ( .A(\myexu/_0017_ ), .Z(\myexu/alu_op [23] ) );
BUF_X1 \myexu/_5326_ ( .A(\src2 [24] ), .Z(\myexu/_2475_ ) );
BUF_X1 \myexu/_5327_ ( .A(\myexu/_0018_ ), .Z(\myexu/alu_op [24] ) );
BUF_X1 \myexu/_5328_ ( .A(\src2 [25] ), .Z(\myexu/_2476_ ) );
BUF_X1 \myexu/_5329_ ( .A(\myexu/_0019_ ), .Z(\myexu/alu_op [25] ) );
BUF_X1 \myexu/_5330_ ( .A(\src2 [26] ), .Z(\myexu/_2477_ ) );
BUF_X1 \myexu/_5331_ ( .A(\myexu/_0020_ ), .Z(\myexu/alu_op [26] ) );
BUF_X1 \myexu/_5332_ ( .A(\src2 [27] ), .Z(\myexu/_2478_ ) );
BUF_X1 \myexu/_5333_ ( .A(\myexu/_0021_ ), .Z(\myexu/alu_op [27] ) );
BUF_X1 \myexu/_5334_ ( .A(\src2 [28] ), .Z(\myexu/_2479_ ) );
BUF_X1 \myexu/_5335_ ( .A(\myexu/_0022_ ), .Z(\myexu/alu_op [28] ) );
BUF_X1 \myexu/_5336_ ( .A(\src2 [29] ), .Z(\myexu/_2480_ ) );
BUF_X1 \myexu/_5337_ ( .A(\myexu/_0023_ ), .Z(\myexu/alu_op [29] ) );
BUF_X1 \myexu/_5338_ ( .A(\src2 [30] ), .Z(\myexu/_2482_ ) );
BUF_X1 \myexu/_5339_ ( .A(\myexu/_0025_ ), .Z(\myexu/alu_op [30] ) );
BUF_X1 \myexu/_5340_ ( .A(\ID_EX_typ [0] ), .Z(\myexu/_2523_ ) );
BUF_X1 \myexu/_5341_ ( .A(\ID_EX_typ [1] ), .Z(\myexu/_2524_ ) );
BUF_X1 \myexu/_5342_ ( .A(\ID_EX_typ [2] ), .Z(\myexu/_2525_ ) );
BUF_X1 \myexu/_5343_ ( .A(\srccs [0] ), .Z(\myexu/_2491_ ) );
BUF_X1 \myexu/_5344_ ( .A(\ID_EX_pc [0] ), .Z(\myexu/_2260_ ) );
BUF_X1 \myexu/_5345_ ( .A(\srccs [1] ), .Z(\myexu/_2502_ ) );
BUF_X1 \myexu/_5346_ ( .A(\ID_EX_pc [1] ), .Z(\myexu/_2271_ ) );
BUF_X1 \myexu/_5347_ ( .A(\srccs [2] ), .Z(\myexu/_2513_ ) );
BUF_X1 \myexu/_5348_ ( .A(\ID_EX_pc [2] ), .Z(\myexu/_2282_ ) );
BUF_X1 \myexu/_5349_ ( .A(\srccs [3] ), .Z(\myexu/_2516_ ) );
BUF_X1 \myexu/_5350_ ( .A(\ID_EX_pc [3] ), .Z(\myexu/_2285_ ) );
BUF_X1 \myexu/_5351_ ( .A(\srccs [4] ), .Z(\myexu/_2517_ ) );
BUF_X1 \myexu/_5352_ ( .A(\ID_EX_pc [4] ), .Z(\myexu/_2286_ ) );
BUF_X1 \myexu/_5353_ ( .A(\srccs [5] ), .Z(\myexu/_2518_ ) );
BUF_X1 \myexu/_5354_ ( .A(\ID_EX_pc [5] ), .Z(\myexu/_2287_ ) );
BUF_X1 \myexu/_5355_ ( .A(\srccs [6] ), .Z(\myexu/_2519_ ) );
BUF_X1 \myexu/_5356_ ( .A(\ID_EX_pc [6] ), .Z(\myexu/_2288_ ) );
BUF_X1 \myexu/_5357_ ( .A(\srccs [7] ), .Z(\myexu/_2520_ ) );
BUF_X1 \myexu/_5358_ ( .A(\ID_EX_pc [7] ), .Z(\myexu/_2289_ ) );
BUF_X1 \myexu/_5359_ ( .A(\srccs [8] ), .Z(\myexu/_2521_ ) );
BUF_X1 \myexu/_5360_ ( .A(\ID_EX_pc [8] ), .Z(\myexu/_2290_ ) );
BUF_X1 \myexu/_5361_ ( .A(\srccs [9] ), .Z(\myexu/_2522_ ) );
BUF_X1 \myexu/_5362_ ( .A(\ID_EX_pc [9] ), .Z(\myexu/_2291_ ) );
BUF_X1 \myexu/_5363_ ( .A(\srccs [10] ), .Z(\myexu/_2492_ ) );
BUF_X1 \myexu/_5364_ ( .A(\ID_EX_pc [10] ), .Z(\myexu/_2261_ ) );
BUF_X1 \myexu/_5365_ ( .A(\srccs [11] ), .Z(\myexu/_2493_ ) );
BUF_X1 \myexu/_5366_ ( .A(\ID_EX_pc [11] ), .Z(\myexu/_2262_ ) );
BUF_X1 \myexu/_5367_ ( .A(\srccs [12] ), .Z(\myexu/_2494_ ) );
BUF_X1 \myexu/_5368_ ( .A(\ID_EX_pc [12] ), .Z(\myexu/_2263_ ) );
BUF_X1 \myexu/_5369_ ( .A(\srccs [13] ), .Z(\myexu/_2495_ ) );
BUF_X1 \myexu/_5370_ ( .A(\ID_EX_pc [13] ), .Z(\myexu/_2264_ ) );
BUF_X1 \myexu/_5371_ ( .A(\srccs [14] ), .Z(\myexu/_2496_ ) );
BUF_X1 \myexu/_5372_ ( .A(\ID_EX_pc [14] ), .Z(\myexu/_2265_ ) );
BUF_X1 \myexu/_5373_ ( .A(\srccs [15] ), .Z(\myexu/_2497_ ) );
BUF_X1 \myexu/_5374_ ( .A(\ID_EX_pc [15] ), .Z(\myexu/_2266_ ) );
BUF_X1 \myexu/_5375_ ( .A(\srccs [16] ), .Z(\myexu/_2498_ ) );
BUF_X1 \myexu/_5376_ ( .A(\ID_EX_pc [16] ), .Z(\myexu/_2267_ ) );
BUF_X1 \myexu/_5377_ ( .A(\srccs [17] ), .Z(\myexu/_2499_ ) );
BUF_X1 \myexu/_5378_ ( .A(\ID_EX_pc [17] ), .Z(\myexu/_2268_ ) );
BUF_X1 \myexu/_5379_ ( .A(\srccs [18] ), .Z(\myexu/_2500_ ) );
BUF_X1 \myexu/_5380_ ( .A(\ID_EX_pc [18] ), .Z(\myexu/_2269_ ) );
BUF_X1 \myexu/_5381_ ( .A(\srccs [19] ), .Z(\myexu/_2501_ ) );
BUF_X1 \myexu/_5382_ ( .A(\ID_EX_pc [19] ), .Z(\myexu/_2270_ ) );
BUF_X1 \myexu/_5383_ ( .A(\srccs [20] ), .Z(\myexu/_2503_ ) );
BUF_X1 \myexu/_5384_ ( .A(\ID_EX_pc [20] ), .Z(\myexu/_2272_ ) );
BUF_X1 \myexu/_5385_ ( .A(\srccs [21] ), .Z(\myexu/_2504_ ) );
BUF_X1 \myexu/_5386_ ( .A(\ID_EX_pc [21] ), .Z(\myexu/_2273_ ) );
BUF_X1 \myexu/_5387_ ( .A(\srccs [22] ), .Z(\myexu/_2505_ ) );
BUF_X1 \myexu/_5388_ ( .A(\ID_EX_pc [22] ), .Z(\myexu/_2274_ ) );
BUF_X1 \myexu/_5389_ ( .A(\srccs [23] ), .Z(\myexu/_2506_ ) );
BUF_X1 \myexu/_5390_ ( .A(\ID_EX_pc [23] ), .Z(\myexu/_2275_ ) );
BUF_X1 \myexu/_5391_ ( .A(\srccs [24] ), .Z(\myexu/_2507_ ) );
BUF_X1 \myexu/_5392_ ( .A(\ID_EX_pc [24] ), .Z(\myexu/_2276_ ) );
BUF_X1 \myexu/_5393_ ( .A(\srccs [25] ), .Z(\myexu/_2508_ ) );
BUF_X1 \myexu/_5394_ ( .A(\ID_EX_pc [25] ), .Z(\myexu/_2277_ ) );
BUF_X1 \myexu/_5395_ ( .A(\srccs [26] ), .Z(\myexu/_2509_ ) );
BUF_X1 \myexu/_5396_ ( .A(\ID_EX_pc [26] ), .Z(\myexu/_2278_ ) );
BUF_X1 \myexu/_5397_ ( .A(\srccs [27] ), .Z(\myexu/_2510_ ) );
BUF_X1 \myexu/_5398_ ( .A(\ID_EX_pc [27] ), .Z(\myexu/_2279_ ) );
BUF_X1 \myexu/_5399_ ( .A(\srccs [28] ), .Z(\myexu/_2511_ ) );
BUF_X1 \myexu/_5400_ ( .A(\ID_EX_pc [28] ), .Z(\myexu/_2280_ ) );
BUF_X1 \myexu/_5401_ ( .A(\srccs [29] ), .Z(\myexu/_2512_ ) );
BUF_X1 \myexu/_5402_ ( .A(\ID_EX_pc [29] ), .Z(\myexu/_2281_ ) );
BUF_X1 \myexu/_5403_ ( .A(\srccs [30] ), .Z(\myexu/_2514_ ) );
BUF_X1 \myexu/_5404_ ( .A(\ID_EX_pc [30] ), .Z(\myexu/_2283_ ) );
BUF_X1 \myexu/_5405_ ( .A(\srccs [31] ), .Z(\myexu/_2515_ ) );
BUF_X1 \myexu/_5406_ ( .A(\ID_EX_pc [31] ), .Z(\myexu/_2284_ ) );
BUF_X1 \myexu/_5407_ ( .A(\ID_EX_csr [0] ), .Z(\myexu/_0243_ ) );
BUF_X1 \myexu/_5408_ ( .A(\ID_EX_csr [1] ), .Z(\myexu/_0246_ ) );
BUF_X1 \myexu/_5409_ ( .A(\ID_EX_csr [2] ), .Z(\myexu/_0247_ ) );
BUF_X1 \myexu/_5410_ ( .A(\ID_EX_csr [3] ), .Z(\myexu/_0248_ ) );
BUF_X1 \myexu/_5411_ ( .A(\ID_EX_csr [4] ), .Z(\myexu/_0249_ ) );
BUF_X1 \myexu/_5412_ ( .A(\ID_EX_csr [5] ), .Z(\myexu/_0250_ ) );
BUF_X1 \myexu/_5413_ ( .A(\ID_EX_csr [6] ), .Z(\myexu/_0251_ ) );
BUF_X1 \myexu/_5414_ ( .A(\ID_EX_csr [7] ), .Z(\myexu/_0252_ ) );
BUF_X1 \myexu/_5415_ ( .A(\ID_EX_csr [8] ), .Z(\myexu/_0253_ ) );
BUF_X1 \myexu/_5416_ ( .A(\ID_EX_csr [9] ), .Z(\myexu/_0254_ ) );
BUF_X1 \myexu/_5417_ ( .A(\ID_EX_csr [10] ), .Z(\myexu/_0244_ ) );
BUF_X1 \myexu/_5418_ ( .A(\ID_EX_csr [11] ), .Z(\myexu/_0245_ ) );
BUF_X1 \myexu/_5419_ ( .A(LSU_arready_set ), .Z(\myexu/_0000_ ) );
BUF_X1 \myexu/_5420_ ( .A(LSU_ready_EXU ), .Z(\myexu/_2361_ ) );
BUF_X1 \myexu/_5421_ ( .A(\EX_LS_flag [0] ), .Z(\myexu/_0292_ ) );
BUF_X1 \myexu/_5422_ ( .A(\EX_LS_flag [1] ), .Z(\myexu/_0293_ ) );
BUF_X1 \myexu/_5423_ ( .A(\EX_LS_flag [2] ), .Z(\myexu/_0294_ ) );
BUF_X1 \myexu/_5424_ ( .A(LSU_awready_set ), .Z(\myexu/_0001_ ) );
BUF_X1 \myexu/_5425_ ( .A(\ID_EX_typ [3] ), .Z(\myexu/_2526_ ) );
BUF_X1 \myexu/_5426_ ( .A(\myexu/alu_out [0] ), .Z(\myexu/_0034_ ) );
BUF_X1 \myexu/_5427_ ( .A(\myexu/alu_out [1] ), .Z(\myexu/_0045_ ) );
BUF_X1 \myexu/_5428_ ( .A(\myexu/alu_out [2] ), .Z(\myexu/_0056_ ) );
BUF_X1 \myexu/_5429_ ( .A(\myexu/alu_out [3] ), .Z(\myexu/_0059_ ) );
BUF_X1 \myexu/_5430_ ( .A(\myexu/alu_out [4] ), .Z(\myexu/_0060_ ) );
BUF_X1 \myexu/_5431_ ( .A(\myexu/alu_out [5] ), .Z(\myexu/_0061_ ) );
BUF_X1 \myexu/_5432_ ( .A(\myexu/alu_out [6] ), .Z(\myexu/_0062_ ) );
BUF_X1 \myexu/_5433_ ( .A(\myexu/alu_out [7] ), .Z(\myexu/_0063_ ) );
BUF_X1 \myexu/_5434_ ( .A(\myexu/alu_out [8] ), .Z(\myexu/_0064_ ) );
BUF_X1 \myexu/_5435_ ( .A(\myexu/alu_out [9] ), .Z(\myexu/_0065_ ) );
BUF_X1 \myexu/_5436_ ( .A(\myexu/alu_out [10] ), .Z(\myexu/_0035_ ) );
BUF_X1 \myexu/_5437_ ( .A(\myexu/alu_out [11] ), .Z(\myexu/_0036_ ) );
BUF_X1 \myexu/_5438_ ( .A(\myexu/alu_out [12] ), .Z(\myexu/_0037_ ) );
BUF_X1 \myexu/_5439_ ( .A(\myexu/alu_out [13] ), .Z(\myexu/_0038_ ) );
BUF_X1 \myexu/_5440_ ( .A(\myexu/alu_out [14] ), .Z(\myexu/_0039_ ) );
BUF_X1 \myexu/_5441_ ( .A(\myexu/alu_out [15] ), .Z(\myexu/_0040_ ) );
BUF_X1 \myexu/_5442_ ( .A(\myexu/alu_out [16] ), .Z(\myexu/_0041_ ) );
BUF_X1 \myexu/_5443_ ( .A(\myexu/alu_out [17] ), .Z(\myexu/_0042_ ) );
BUF_X1 \myexu/_5444_ ( .A(\myexu/alu_out [18] ), .Z(\myexu/_0043_ ) );
BUF_X1 \myexu/_5445_ ( .A(\myexu/alu_out [19] ), .Z(\myexu/_0044_ ) );
BUF_X1 \myexu/_5446_ ( .A(\myexu/alu_out [20] ), .Z(\myexu/_0046_ ) );
BUF_X1 \myexu/_5447_ ( .A(\myexu/alu_out [21] ), .Z(\myexu/_0047_ ) );
BUF_X1 \myexu/_5448_ ( .A(\myexu/alu_out [22] ), .Z(\myexu/_0048_ ) );
BUF_X1 \myexu/_5449_ ( .A(\myexu/alu_out [23] ), .Z(\myexu/_0049_ ) );
BUF_X1 \myexu/_5450_ ( .A(\myexu/alu_out [24] ), .Z(\myexu/_0050_ ) );
BUF_X1 \myexu/_5451_ ( .A(\myexu/alu_out [25] ), .Z(\myexu/_0051_ ) );
BUF_X1 \myexu/_5452_ ( .A(\myexu/alu_out [26] ), .Z(\myexu/_0052_ ) );
BUF_X1 \myexu/_5453_ ( .A(\myexu/alu_out [27] ), .Z(\myexu/_0053_ ) );
BUF_X1 \myexu/_5454_ ( .A(\myexu/alu_out [28] ), .Z(\myexu/_0054_ ) );
BUF_X1 \myexu/_5455_ ( .A(\myexu/alu_out [29] ), .Z(\myexu/_0055_ ) );
BUF_X1 \myexu/_5456_ ( .A(\myexu/alu_out [30] ), .Z(\myexu/_0057_ ) );
BUF_X1 \myexu/_5457_ ( .A(\myexu/alu_out [31] ), .Z(\myexu/_0058_ ) );
BUF_X1 \myexu/_5458_ ( .A(check_quest ), .Z(\myexu/_0242_ ) );
BUF_X1 \myexu/_5459_ ( .A(check_assert ), .Z(\myexu/_0241_ ) );
BUF_X1 \myexu/_5460_ ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(\myexu/_0255_ ) );
BUF_X1 \myexu/_5461_ ( .A(\myexu/_0066_ ), .Z(\myexu/_2712_ ) );
BUF_X1 \myexu/_5462_ ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(\myexu/_0266_ ) );
BUF_X1 \myexu/_5463_ ( .A(\myexu/_0067_ ), .Z(\myexu/_2713_ ) );
BUF_X1 \myexu/_5464_ ( .A(\EX_LS_dest_csreg_mem [2] ), .Z(\myexu/_0277_ ) );
BUF_X1 \myexu/_5465_ ( .A(\myexu/_0068_ ), .Z(\myexu/_2714_ ) );
BUF_X1 \myexu/_5466_ ( .A(\EX_LS_dest_csreg_mem [3] ), .Z(\myexu/_0280_ ) );
BUF_X1 \myexu/_5467_ ( .A(\myexu/_0069_ ), .Z(\myexu/_2715_ ) );
BUF_X1 \myexu/_5468_ ( .A(\EX_LS_dest_csreg_mem [4] ), .Z(\myexu/_0281_ ) );
BUF_X1 \myexu/_5469_ ( .A(\myexu/_0070_ ), .Z(\myexu/_2716_ ) );
BUF_X1 \myexu/_5470_ ( .A(\EX_LS_dest_csreg_mem [5] ), .Z(\myexu/_0282_ ) );
BUF_X1 \myexu/_5471_ ( .A(\myexu/_0071_ ), .Z(\myexu/_2717_ ) );
BUF_X1 \myexu/_5472_ ( .A(\EX_LS_dest_csreg_mem [6] ), .Z(\myexu/_0283_ ) );
BUF_X1 \myexu/_5473_ ( .A(\myexu/_0072_ ), .Z(\myexu/_2718_ ) );
BUF_X1 \myexu/_5474_ ( .A(\EX_LS_dest_csreg_mem [7] ), .Z(\myexu/_0284_ ) );
BUF_X1 \myexu/_5475_ ( .A(\myexu/_0073_ ), .Z(\myexu/_2719_ ) );
BUF_X1 \myexu/_5476_ ( .A(\EX_LS_dest_csreg_mem [8] ), .Z(\myexu/_0285_ ) );
BUF_X1 \myexu/_5477_ ( .A(\myexu/_0074_ ), .Z(\myexu/_2720_ ) );
BUF_X1 \myexu/_5478_ ( .A(\EX_LS_dest_csreg_mem [9] ), .Z(\myexu/_0286_ ) );
BUF_X1 \myexu/_5479_ ( .A(\myexu/_0075_ ), .Z(\myexu/_2721_ ) );
BUF_X1 \myexu/_5480_ ( .A(\EX_LS_dest_csreg_mem [10] ), .Z(\myexu/_0256_ ) );
BUF_X1 \myexu/_5481_ ( .A(\myexu/_0076_ ), .Z(\myexu/_2722_ ) );
BUF_X1 \myexu/_5482_ ( .A(\EX_LS_dest_csreg_mem [11] ), .Z(\myexu/_0257_ ) );
BUF_X1 \myexu/_5483_ ( .A(\myexu/_0077_ ), .Z(\myexu/_2723_ ) );
BUF_X1 \myexu/_5484_ ( .A(\EX_LS_result_csreg_mem [0] ), .Z(\myexu/_2362_ ) );
BUF_X1 \myexu/_5485_ ( .A(\myexu/_0078_ ), .Z(\myexu/_2724_ ) );
BUF_X1 \myexu/_5486_ ( .A(\EX_LS_result_csreg_mem [1] ), .Z(\myexu/_2373_ ) );
BUF_X1 \myexu/_5487_ ( .A(\myexu/_0079_ ), .Z(\myexu/_2725_ ) );
BUF_X1 \myexu/_5488_ ( .A(\EX_LS_result_csreg_mem [2] ), .Z(\myexu/_2384_ ) );
BUF_X1 \myexu/_5489_ ( .A(\myexu/_0080_ ), .Z(\myexu/_2726_ ) );
BUF_X1 \myexu/_5490_ ( .A(\EX_LS_result_csreg_mem [3] ), .Z(\myexu/_2387_ ) );
BUF_X1 \myexu/_5491_ ( .A(\myexu/_0081_ ), .Z(\myexu/_2727_ ) );
BUF_X1 \myexu/_5492_ ( .A(\EX_LS_result_csreg_mem [4] ), .Z(\myexu/_2388_ ) );
BUF_X1 \myexu/_5493_ ( .A(\myexu/_0082_ ), .Z(\myexu/_2728_ ) );
BUF_X1 \myexu/_5494_ ( .A(\EX_LS_result_csreg_mem [5] ), .Z(\myexu/_2389_ ) );
BUF_X1 \myexu/_5495_ ( .A(\myexu/_0083_ ), .Z(\myexu/_2729_ ) );
BUF_X1 \myexu/_5496_ ( .A(\EX_LS_result_csreg_mem [6] ), .Z(\myexu/_2390_ ) );
BUF_X1 \myexu/_5497_ ( .A(\myexu/_0084_ ), .Z(\myexu/_2730_ ) );
BUF_X1 \myexu/_5498_ ( .A(\EX_LS_result_csreg_mem [7] ), .Z(\myexu/_2391_ ) );
BUF_X1 \myexu/_5499_ ( .A(\myexu/_0085_ ), .Z(\myexu/_2731_ ) );
BUF_X1 \myexu/_5500_ ( .A(\EX_LS_result_csreg_mem [8] ), .Z(\myexu/_2392_ ) );
BUF_X1 \myexu/_5501_ ( .A(\myexu/_0086_ ), .Z(\myexu/_2732_ ) );
BUF_X1 \myexu/_5502_ ( .A(\EX_LS_result_csreg_mem [9] ), .Z(\myexu/_2393_ ) );
BUF_X1 \myexu/_5503_ ( .A(\myexu/_0087_ ), .Z(\myexu/_2733_ ) );
BUF_X1 \myexu/_5504_ ( .A(\EX_LS_result_csreg_mem [10] ), .Z(\myexu/_2363_ ) );
BUF_X1 \myexu/_5505_ ( .A(\myexu/_0088_ ), .Z(\myexu/_2734_ ) );
BUF_X1 \myexu/_5506_ ( .A(\EX_LS_result_csreg_mem [11] ), .Z(\myexu/_2364_ ) );
BUF_X1 \myexu/_5507_ ( .A(\myexu/_0089_ ), .Z(\myexu/_2735_ ) );
BUF_X1 \myexu/_5508_ ( .A(\EX_LS_result_csreg_mem [12] ), .Z(\myexu/_2365_ ) );
BUF_X1 \myexu/_5509_ ( .A(\myexu/_0090_ ), .Z(\myexu/_2736_ ) );
BUF_X1 \myexu/_5510_ ( .A(\EX_LS_result_csreg_mem [13] ), .Z(\myexu/_2366_ ) );
BUF_X1 \myexu/_5511_ ( .A(\myexu/_0091_ ), .Z(\myexu/_2737_ ) );
BUF_X1 \myexu/_5512_ ( .A(\EX_LS_result_csreg_mem [14] ), .Z(\myexu/_2367_ ) );
BUF_X1 \myexu/_5513_ ( .A(\myexu/_0092_ ), .Z(\myexu/_2738_ ) );
BUF_X1 \myexu/_5514_ ( .A(\EX_LS_result_csreg_mem [15] ), .Z(\myexu/_2368_ ) );
BUF_X1 \myexu/_5515_ ( .A(\myexu/_0093_ ), .Z(\myexu/_2739_ ) );
BUF_X1 \myexu/_5516_ ( .A(\EX_LS_result_csreg_mem [16] ), .Z(\myexu/_2369_ ) );
BUF_X1 \myexu/_5517_ ( .A(\myexu/_0094_ ), .Z(\myexu/_2740_ ) );
BUF_X1 \myexu/_5518_ ( .A(\EX_LS_result_csreg_mem [17] ), .Z(\myexu/_2370_ ) );
BUF_X1 \myexu/_5519_ ( .A(\myexu/_0095_ ), .Z(\myexu/_2741_ ) );
BUF_X1 \myexu/_5520_ ( .A(\EX_LS_result_csreg_mem [18] ), .Z(\myexu/_2371_ ) );
BUF_X1 \myexu/_5521_ ( .A(\myexu/_0096_ ), .Z(\myexu/_2742_ ) );
BUF_X1 \myexu/_5522_ ( .A(\EX_LS_result_csreg_mem [19] ), .Z(\myexu/_2372_ ) );
BUF_X1 \myexu/_5523_ ( .A(\myexu/_0097_ ), .Z(\myexu/_2743_ ) );
BUF_X1 \myexu/_5524_ ( .A(\EX_LS_result_csreg_mem [20] ), .Z(\myexu/_2374_ ) );
BUF_X1 \myexu/_5525_ ( .A(\myexu/_0098_ ), .Z(\myexu/_2744_ ) );
BUF_X1 \myexu/_5526_ ( .A(\EX_LS_result_csreg_mem [21] ), .Z(\myexu/_2375_ ) );
BUF_X1 \myexu/_5527_ ( .A(\myexu/_0099_ ), .Z(\myexu/_2745_ ) );
BUF_X1 \myexu/_5528_ ( .A(\EX_LS_result_csreg_mem [22] ), .Z(\myexu/_2376_ ) );
BUF_X1 \myexu/_5529_ ( .A(\myexu/_0100_ ), .Z(\myexu/_2746_ ) );
BUF_X1 \myexu/_5530_ ( .A(\EX_LS_result_csreg_mem [23] ), .Z(\myexu/_2377_ ) );
BUF_X1 \myexu/_5531_ ( .A(\myexu/_0101_ ), .Z(\myexu/_2747_ ) );
BUF_X1 \myexu/_5532_ ( .A(\EX_LS_result_csreg_mem [24] ), .Z(\myexu/_2378_ ) );
BUF_X1 \myexu/_5533_ ( .A(\myexu/_0102_ ), .Z(\myexu/_2748_ ) );
BUF_X1 \myexu/_5534_ ( .A(\EX_LS_result_csreg_mem [25] ), .Z(\myexu/_2379_ ) );
BUF_X1 \myexu/_5535_ ( .A(\myexu/_0103_ ), .Z(\myexu/_2749_ ) );
BUF_X1 \myexu/_5536_ ( .A(\EX_LS_result_csreg_mem [26] ), .Z(\myexu/_2380_ ) );
BUF_X1 \myexu/_5537_ ( .A(\myexu/_0104_ ), .Z(\myexu/_2750_ ) );
BUF_X1 \myexu/_5538_ ( .A(\EX_LS_result_csreg_mem [27] ), .Z(\myexu/_2381_ ) );
BUF_X1 \myexu/_5539_ ( .A(\myexu/_0105_ ), .Z(\myexu/_2751_ ) );
BUF_X1 \myexu/_5540_ ( .A(\EX_LS_result_csreg_mem [28] ), .Z(\myexu/_2382_ ) );
BUF_X1 \myexu/_5541_ ( .A(\myexu/_0106_ ), .Z(\myexu/_2752_ ) );
BUF_X1 \myexu/_5542_ ( .A(\EX_LS_result_csreg_mem [29] ), .Z(\myexu/_2383_ ) );
BUF_X1 \myexu/_5543_ ( .A(\myexu/_0107_ ), .Z(\myexu/_2753_ ) );
BUF_X1 \myexu/_5544_ ( .A(\EX_LS_result_csreg_mem [30] ), .Z(\myexu/_2385_ ) );
BUF_X1 \myexu/_5545_ ( .A(\myexu/_0108_ ), .Z(\myexu/_2754_ ) );
BUF_X1 \myexu/_5546_ ( .A(\EX_LS_result_csreg_mem [31] ), .Z(\myexu/_2386_ ) );
BUF_X1 \myexu/_5547_ ( .A(\myexu/_0109_ ), .Z(\myexu/_2755_ ) );
BUF_X1 \myexu/_5548_ ( .A(\pc_jump [0] ), .Z(\myexu/_2292_ ) );
BUF_X1 \myexu/_5549_ ( .A(\pc_jump [1] ), .Z(\myexu/_2303_ ) );
BUF_X1 \myexu/_5550_ ( .A(\pc_jump [2] ), .Z(\myexu/_2314_ ) );
BUF_X1 \myexu/_5551_ ( .A(\pc_jump [3] ), .Z(\myexu/_2317_ ) );
BUF_X1 \myexu/_5552_ ( .A(\pc_jump [4] ), .Z(\myexu/_2318_ ) );
BUF_X1 \myexu/_5553_ ( .A(\pc_jump [5] ), .Z(\myexu/_2319_ ) );
BUF_X1 \myexu/_5554_ ( .A(\pc_jump [6] ), .Z(\myexu/_2320_ ) );
BUF_X1 \myexu/_5555_ ( .A(\pc_jump [7] ), .Z(\myexu/_2321_ ) );
BUF_X1 \myexu/_5556_ ( .A(\pc_jump [8] ), .Z(\myexu/_2322_ ) );
BUF_X1 \myexu/_5557_ ( .A(\pc_jump [9] ), .Z(\myexu/_2323_ ) );
BUF_X1 \myexu/_5558_ ( .A(\pc_jump [10] ), .Z(\myexu/_2293_ ) );
BUF_X1 \myexu/_5559_ ( .A(\pc_jump [11] ), .Z(\myexu/_2294_ ) );
BUF_X1 \myexu/_5560_ ( .A(\pc_jump [12] ), .Z(\myexu/_2295_ ) );
BUF_X1 \myexu/_5561_ ( .A(\pc_jump [13] ), .Z(\myexu/_2296_ ) );
BUF_X1 \myexu/_5562_ ( .A(\pc_jump [14] ), .Z(\myexu/_2297_ ) );
BUF_X1 \myexu/_5563_ ( .A(\pc_jump [15] ), .Z(\myexu/_2298_ ) );
BUF_X1 \myexu/_5564_ ( .A(\pc_jump [16] ), .Z(\myexu/_2299_ ) );
BUF_X1 \myexu/_5565_ ( .A(\pc_jump [17] ), .Z(\myexu/_2300_ ) );
BUF_X1 \myexu/_5566_ ( .A(\pc_jump [18] ), .Z(\myexu/_2301_ ) );
BUF_X1 \myexu/_5567_ ( .A(\pc_jump [19] ), .Z(\myexu/_2302_ ) );
BUF_X1 \myexu/_5568_ ( .A(\pc_jump [20] ), .Z(\myexu/_2304_ ) );
BUF_X1 \myexu/_5569_ ( .A(\pc_jump [21] ), .Z(\myexu/_2305_ ) );
BUF_X1 \myexu/_5570_ ( .A(\pc_jump [22] ), .Z(\myexu/_2306_ ) );
BUF_X1 \myexu/_5571_ ( .A(\pc_jump [23] ), .Z(\myexu/_2307_ ) );
BUF_X1 \myexu/_5572_ ( .A(\pc_jump [24] ), .Z(\myexu/_2308_ ) );
BUF_X1 \myexu/_5573_ ( .A(\pc_jump [25] ), .Z(\myexu/_2309_ ) );
BUF_X1 \myexu/_5574_ ( .A(\pc_jump [26] ), .Z(\myexu/_2310_ ) );
BUF_X1 \myexu/_5575_ ( .A(\pc_jump [27] ), .Z(\myexu/_2311_ ) );
BUF_X1 \myexu/_5576_ ( .A(\pc_jump [28] ), .Z(\myexu/_2312_ ) );
BUF_X1 \myexu/_5577_ ( .A(\pc_jump [29] ), .Z(\myexu/_2313_ ) );
BUF_X1 \myexu/_5578_ ( .A(\pc_jump [30] ), .Z(\myexu/_2315_ ) );
BUF_X1 \myexu/_5579_ ( .A(\pc_jump [31] ), .Z(\myexu/_2316_ ) );
BUF_X1 \myexu/_5580_ ( .A(\EX_LS_pc [0] ), .Z(\myexu/_2324_ ) );
BUF_X1 \myexu/_5581_ ( .A(\EX_LS_pc [1] ), .Z(\myexu/_2335_ ) );
BUF_X1 \myexu/_5582_ ( .A(\EX_LS_pc [2] ), .Z(\myexu/_2346_ ) );
BUF_X1 \myexu/_5583_ ( .A(\EX_LS_pc [3] ), .Z(\myexu/_2349_ ) );
BUF_X1 \myexu/_5584_ ( .A(\EX_LS_pc [4] ), .Z(\myexu/_2350_ ) );
BUF_X1 \myexu/_5585_ ( .A(\EX_LS_pc [5] ), .Z(\myexu/_2351_ ) );
BUF_X1 \myexu/_5586_ ( .A(\EX_LS_pc [6] ), .Z(\myexu/_2352_ ) );
BUF_X1 \myexu/_5587_ ( .A(\EX_LS_pc [7] ), .Z(\myexu/_2353_ ) );
BUF_X1 \myexu/_5588_ ( .A(\EX_LS_pc [8] ), .Z(\myexu/_2354_ ) );
BUF_X1 \myexu/_5589_ ( .A(\EX_LS_pc [9] ), .Z(\myexu/_2355_ ) );
BUF_X1 \myexu/_5590_ ( .A(\EX_LS_pc [10] ), .Z(\myexu/_2325_ ) );
BUF_X1 \myexu/_5591_ ( .A(\EX_LS_pc [11] ), .Z(\myexu/_2326_ ) );
BUF_X1 \myexu/_5592_ ( .A(\EX_LS_pc [12] ), .Z(\myexu/_2327_ ) );
BUF_X1 \myexu/_5593_ ( .A(\EX_LS_pc [13] ), .Z(\myexu/_2328_ ) );
BUF_X1 \myexu/_5594_ ( .A(\EX_LS_pc [14] ), .Z(\myexu/_2329_ ) );
BUF_X1 \myexu/_5595_ ( .A(\EX_LS_pc [15] ), .Z(\myexu/_2330_ ) );
BUF_X1 \myexu/_5596_ ( .A(\EX_LS_pc [16] ), .Z(\myexu/_2331_ ) );
BUF_X1 \myexu/_5597_ ( .A(\EX_LS_pc [17] ), .Z(\myexu/_2332_ ) );
BUF_X1 \myexu/_5598_ ( .A(\EX_LS_pc [18] ), .Z(\myexu/_2333_ ) );
BUF_X1 \myexu/_5599_ ( .A(\EX_LS_pc [19] ), .Z(\myexu/_2334_ ) );
BUF_X1 \myexu/_5600_ ( .A(\EX_LS_pc [20] ), .Z(\myexu/_2336_ ) );
BUF_X1 \myexu/_5601_ ( .A(\EX_LS_pc [21] ), .Z(\myexu/_2337_ ) );
BUF_X1 \myexu/_5602_ ( .A(\EX_LS_pc [22] ), .Z(\myexu/_2338_ ) );
BUF_X1 \myexu/_5603_ ( .A(\EX_LS_pc [23] ), .Z(\myexu/_2339_ ) );
BUF_X1 \myexu/_5604_ ( .A(\EX_LS_pc [24] ), .Z(\myexu/_2340_ ) );
BUF_X1 \myexu/_5605_ ( .A(\EX_LS_pc [25] ), .Z(\myexu/_2341_ ) );
BUF_X1 \myexu/_5606_ ( .A(\EX_LS_pc [26] ), .Z(\myexu/_2342_ ) );
BUF_X1 \myexu/_5607_ ( .A(\EX_LS_pc [27] ), .Z(\myexu/_2343_ ) );
BUF_X1 \myexu/_5608_ ( .A(\EX_LS_pc [28] ), .Z(\myexu/_2344_ ) );
BUF_X1 \myexu/_5609_ ( .A(\EX_LS_pc [29] ), .Z(\myexu/_2345_ ) );
BUF_X1 \myexu/_5610_ ( .A(\EX_LS_pc [30] ), .Z(\myexu/_2347_ ) );
BUF_X1 \myexu/_5611_ ( .A(\EX_LS_pc [31] ), .Z(\myexu/_2348_ ) );
BUF_X1 \myexu/_5612_ ( .A(\EX_LS_typ [0] ), .Z(\myexu/_2531_ ) );
BUF_X1 \myexu/_5613_ ( .A(\EX_LS_typ [1] ), .Z(\myexu/_2532_ ) );
BUF_X1 \myexu/_5614_ ( .A(\EX_LS_typ [2] ), .Z(\myexu/_2533_ ) );
BUF_X1 \myexu/_5615_ ( .A(\EX_LS_typ [3] ), .Z(\myexu/_2534_ ) );
BUF_X1 \myexu/_5616_ ( .A(\EX_LS_typ [4] ), .Z(\myexu/_2535_ ) );
BUF_X1 \myexu/_5617_ ( .A(\EX_LS_dest_reg [0] ), .Z(\myexu/_0287_ ) );
BUF_X1 \myexu/_5618_ ( .A(\ID_EX_rd [0] ), .Z(\myexu/_2356_ ) );
BUF_X1 \myexu/_5619_ ( .A(\EX_LS_dest_reg [1] ), .Z(\myexu/_0288_ ) );
BUF_X1 \myexu/_5620_ ( .A(\ID_EX_rd [1] ), .Z(\myexu/_2357_ ) );
BUF_X1 \myexu/_5621_ ( .A(\EX_LS_dest_reg [2] ), .Z(\myexu/_0289_ ) );
BUF_X1 \myexu/_5622_ ( .A(\ID_EX_rd [2] ), .Z(\myexu/_2358_ ) );
BUF_X1 \myexu/_5623_ ( .A(\EX_LS_dest_reg [3] ), .Z(\myexu/_0290_ ) );
BUF_X1 \myexu/_5624_ ( .A(\ID_EX_rd [3] ), .Z(\myexu/_2359_ ) );
BUF_X1 \myexu/_5625_ ( .A(\EX_LS_dest_reg [4] ), .Z(\myexu/_0291_ ) );
BUF_X1 \myexu/_5626_ ( .A(\ID_EX_rd [4] ), .Z(\myexu/_2360_ ) );
BUF_X1 \myexu/_5627_ ( .A(\EX_LS_dest_csreg_mem [12] ), .Z(\myexu/_0258_ ) );
BUF_X1 \myexu/_5628_ ( .A(\myexu/_0189_ ), .Z(\myexu/_2835_ ) );
BUF_X1 \myexu/_5629_ ( .A(\EX_LS_dest_csreg_mem [13] ), .Z(\myexu/_0259_ ) );
BUF_X1 \myexu/_5630_ ( .A(\myexu/_0190_ ), .Z(\myexu/_2836_ ) );
BUF_X1 \myexu/_5631_ ( .A(\EX_LS_dest_csreg_mem [14] ), .Z(\myexu/_0260_ ) );
BUF_X1 \myexu/_5632_ ( .A(\myexu/_0191_ ), .Z(\myexu/_2837_ ) );
BUF_X1 \myexu/_5633_ ( .A(\EX_LS_dest_csreg_mem [15] ), .Z(\myexu/_0261_ ) );
BUF_X1 \myexu/_5634_ ( .A(\myexu/_0192_ ), .Z(\myexu/_2838_ ) );
BUF_X1 \myexu/_5635_ ( .A(\EX_LS_dest_csreg_mem [16] ), .Z(\myexu/_0262_ ) );
BUF_X1 \myexu/_5636_ ( .A(\myexu/_0193_ ), .Z(\myexu/_2839_ ) );
BUF_X1 \myexu/_5637_ ( .A(\EX_LS_dest_csreg_mem [17] ), .Z(\myexu/_0263_ ) );
BUF_X1 \myexu/_5638_ ( .A(\myexu/_0194_ ), .Z(\myexu/_2840_ ) );
BUF_X1 \myexu/_5639_ ( .A(\EX_LS_dest_csreg_mem [18] ), .Z(\myexu/_0264_ ) );
BUF_X1 \myexu/_5640_ ( .A(\myexu/_0195_ ), .Z(\myexu/_2841_ ) );
BUF_X1 \myexu/_5641_ ( .A(\EX_LS_dest_csreg_mem [19] ), .Z(\myexu/_0265_ ) );
BUF_X1 \myexu/_5642_ ( .A(\myexu/_0196_ ), .Z(\myexu/_2842_ ) );
BUF_X1 \myexu/_5643_ ( .A(\EX_LS_dest_csreg_mem [20] ), .Z(\myexu/_0267_ ) );
BUF_X1 \myexu/_5644_ ( .A(\myexu/_0197_ ), .Z(\myexu/_2843_ ) );
BUF_X1 \myexu/_5645_ ( .A(\EX_LS_dest_csreg_mem [21] ), .Z(\myexu/_0268_ ) );
BUF_X1 \myexu/_5646_ ( .A(\myexu/_0198_ ), .Z(\myexu/_2844_ ) );
BUF_X1 \myexu/_5647_ ( .A(\EX_LS_dest_csreg_mem [22] ), .Z(\myexu/_0269_ ) );
BUF_X1 \myexu/_5648_ ( .A(\myexu/_0199_ ), .Z(\myexu/_2845_ ) );
BUF_X1 \myexu/_5649_ ( .A(\EX_LS_dest_csreg_mem [23] ), .Z(\myexu/_0270_ ) );
BUF_X1 \myexu/_5650_ ( .A(\myexu/_0200_ ), .Z(\myexu/_2846_ ) );
BUF_X1 \myexu/_5651_ ( .A(\EX_LS_dest_csreg_mem [24] ), .Z(\myexu/_0271_ ) );
BUF_X1 \myexu/_5652_ ( .A(\myexu/_0201_ ), .Z(\myexu/_2847_ ) );
BUF_X1 \myexu/_5653_ ( .A(\EX_LS_dest_csreg_mem [25] ), .Z(\myexu/_0272_ ) );
BUF_X1 \myexu/_5654_ ( .A(\myexu/_0202_ ), .Z(\myexu/_2848_ ) );
BUF_X1 \myexu/_5655_ ( .A(\EX_LS_dest_csreg_mem [26] ), .Z(\myexu/_0273_ ) );
BUF_X1 \myexu/_5656_ ( .A(\myexu/_0203_ ), .Z(\myexu/_2849_ ) );
BUF_X1 \myexu/_5657_ ( .A(\EX_LS_dest_csreg_mem [27] ), .Z(\myexu/_0274_ ) );
BUF_X1 \myexu/_5658_ ( .A(\myexu/_0204_ ), .Z(\myexu/_2850_ ) );
BUF_X1 \myexu/_5659_ ( .A(\EX_LS_dest_csreg_mem [28] ), .Z(\myexu/_0275_ ) );
BUF_X1 \myexu/_5660_ ( .A(\myexu/_0205_ ), .Z(\myexu/_2851_ ) );
BUF_X1 \myexu/_5661_ ( .A(\EX_LS_dest_csreg_mem [29] ), .Z(\myexu/_0276_ ) );
BUF_X1 \myexu/_5662_ ( .A(\myexu/_0206_ ), .Z(\myexu/_2852_ ) );
BUF_X1 \myexu/_5663_ ( .A(\EX_LS_dest_csreg_mem [30] ), .Z(\myexu/_0278_ ) );
BUF_X1 \myexu/_5664_ ( .A(\myexu/_0207_ ), .Z(\myexu/_2853_ ) );
BUF_X1 \myexu/_5665_ ( .A(\EX_LS_dest_csreg_mem [31] ), .Z(\myexu/_0279_ ) );
BUF_X1 \myexu/_5666_ ( .A(\myexu/_0208_ ), .Z(\myexu/_2854_ ) );
BUF_X1 \myexu/_5667_ ( .A(\EX_LS_result_reg [0] ), .Z(\myexu/_2394_ ) );
BUF_X1 \myexu/_5668_ ( .A(\myexu/_0209_ ), .Z(\myexu/_2855_ ) );
BUF_X1 \myexu/_5669_ ( .A(\EX_LS_result_reg [1] ), .Z(\myexu/_2405_ ) );
BUF_X1 \myexu/_5670_ ( .A(\myexu/_0210_ ), .Z(\myexu/_2856_ ) );
BUF_X1 \myexu/_5671_ ( .A(\EX_LS_result_reg [2] ), .Z(\myexu/_2416_ ) );
BUF_X1 \myexu/_5672_ ( .A(\myexu/_0211_ ), .Z(\myexu/_2857_ ) );
BUF_X1 \myexu/_5673_ ( .A(\EX_LS_result_reg [3] ), .Z(\myexu/_2419_ ) );
BUF_X1 \myexu/_5674_ ( .A(\myexu/_0212_ ), .Z(\myexu/_2858_ ) );
BUF_X1 \myexu/_5675_ ( .A(\EX_LS_result_reg [4] ), .Z(\myexu/_2420_ ) );
BUF_X1 \myexu/_5676_ ( .A(\myexu/_0213_ ), .Z(\myexu/_2859_ ) );
BUF_X1 \myexu/_5677_ ( .A(\EX_LS_result_reg [5] ), .Z(\myexu/_2421_ ) );
BUF_X1 \myexu/_5678_ ( .A(\myexu/_0214_ ), .Z(\myexu/_2860_ ) );
BUF_X1 \myexu/_5679_ ( .A(\EX_LS_result_reg [6] ), .Z(\myexu/_2422_ ) );
BUF_X1 \myexu/_5680_ ( .A(\myexu/_0215_ ), .Z(\myexu/_2861_ ) );
BUF_X1 \myexu/_5681_ ( .A(\EX_LS_result_reg [7] ), .Z(\myexu/_2423_ ) );
BUF_X1 \myexu/_5682_ ( .A(\myexu/_0216_ ), .Z(\myexu/_2862_ ) );
BUF_X1 \myexu/_5683_ ( .A(\EX_LS_result_reg [8] ), .Z(\myexu/_2424_ ) );
BUF_X1 \myexu/_5684_ ( .A(\myexu/_0217_ ), .Z(\myexu/_2863_ ) );
BUF_X1 \myexu/_5685_ ( .A(\EX_LS_result_reg [9] ), .Z(\myexu/_2425_ ) );
BUF_X1 \myexu/_5686_ ( .A(\myexu/_0218_ ), .Z(\myexu/_2864_ ) );
BUF_X1 \myexu/_5687_ ( .A(\EX_LS_result_reg [10] ), .Z(\myexu/_2395_ ) );
BUF_X1 \myexu/_5688_ ( .A(\myexu/_0219_ ), .Z(\myexu/_2865_ ) );
BUF_X1 \myexu/_5689_ ( .A(\EX_LS_result_reg [11] ), .Z(\myexu/_2396_ ) );
BUF_X1 \myexu/_5690_ ( .A(\myexu/_0220_ ), .Z(\myexu/_2866_ ) );
BUF_X1 \myexu/_5691_ ( .A(\EX_LS_result_reg [12] ), .Z(\myexu/_2397_ ) );
BUF_X1 \myexu/_5692_ ( .A(\myexu/_0221_ ), .Z(\myexu/_2867_ ) );
BUF_X1 \myexu/_5693_ ( .A(\EX_LS_result_reg [13] ), .Z(\myexu/_2398_ ) );
BUF_X1 \myexu/_5694_ ( .A(\myexu/_0222_ ), .Z(\myexu/_2868_ ) );
BUF_X1 \myexu/_5695_ ( .A(\EX_LS_result_reg [14] ), .Z(\myexu/_2399_ ) );
BUF_X1 \myexu/_5696_ ( .A(\myexu/_0223_ ), .Z(\myexu/_2869_ ) );
BUF_X1 \myexu/_5697_ ( .A(\EX_LS_result_reg [15] ), .Z(\myexu/_2400_ ) );
BUF_X1 \myexu/_5698_ ( .A(\myexu/_0224_ ), .Z(\myexu/_2870_ ) );
BUF_X1 \myexu/_5699_ ( .A(\EX_LS_result_reg [16] ), .Z(\myexu/_2401_ ) );
BUF_X1 \myexu/_5700_ ( .A(\myexu/_0225_ ), .Z(\myexu/_2871_ ) );
BUF_X1 \myexu/_5701_ ( .A(\EX_LS_result_reg [17] ), .Z(\myexu/_2402_ ) );
BUF_X1 \myexu/_5702_ ( .A(\myexu/_0226_ ), .Z(\myexu/_2872_ ) );
BUF_X1 \myexu/_5703_ ( .A(\EX_LS_result_reg [18] ), .Z(\myexu/_2403_ ) );
BUF_X1 \myexu/_5704_ ( .A(\myexu/_0227_ ), .Z(\myexu/_2873_ ) );
BUF_X1 \myexu/_5705_ ( .A(\EX_LS_result_reg [19] ), .Z(\myexu/_2404_ ) );
BUF_X1 \myexu/_5706_ ( .A(\myexu/_0228_ ), .Z(\myexu/_2874_ ) );
BUF_X1 \myexu/_5707_ ( .A(\EX_LS_result_reg [20] ), .Z(\myexu/_2406_ ) );
BUF_X1 \myexu/_5708_ ( .A(\myexu/_0229_ ), .Z(\myexu/_2875_ ) );
BUF_X1 \myexu/_5709_ ( .A(\EX_LS_result_reg [21] ), .Z(\myexu/_2407_ ) );
BUF_X1 \myexu/_5710_ ( .A(\myexu/_0230_ ), .Z(\myexu/_2876_ ) );
BUF_X1 \myexu/_5711_ ( .A(\EX_LS_result_reg [22] ), .Z(\myexu/_2408_ ) );
BUF_X1 \myexu/_5712_ ( .A(\myexu/_0231_ ), .Z(\myexu/_2877_ ) );
BUF_X1 \myexu/_5713_ ( .A(\EX_LS_result_reg [23] ), .Z(\myexu/_2409_ ) );
BUF_X1 \myexu/_5714_ ( .A(\myexu/_0232_ ), .Z(\myexu/_2878_ ) );
BUF_X1 \myexu/_5715_ ( .A(\EX_LS_result_reg [24] ), .Z(\myexu/_2410_ ) );
BUF_X1 \myexu/_5716_ ( .A(\myexu/_0233_ ), .Z(\myexu/_2879_ ) );
BUF_X1 \myexu/_5717_ ( .A(\EX_LS_result_reg [25] ), .Z(\myexu/_2411_ ) );
BUF_X1 \myexu/_5718_ ( .A(\myexu/_0234_ ), .Z(\myexu/_2880_ ) );
BUF_X1 \myexu/_5719_ ( .A(\EX_LS_result_reg [26] ), .Z(\myexu/_2412_ ) );
BUF_X1 \myexu/_5720_ ( .A(\myexu/_0235_ ), .Z(\myexu/_2881_ ) );
BUF_X1 \myexu/_5721_ ( .A(\EX_LS_result_reg [27] ), .Z(\myexu/_2413_ ) );
BUF_X1 \myexu/_5722_ ( .A(\myexu/_0236_ ), .Z(\myexu/_2882_ ) );
BUF_X1 \myexu/_5723_ ( .A(\EX_LS_result_reg [28] ), .Z(\myexu/_2414_ ) );
BUF_X1 \myexu/_5724_ ( .A(\myexu/_0237_ ), .Z(\myexu/_2883_ ) );
BUF_X1 \myexu/_5725_ ( .A(\EX_LS_result_reg [29] ), .Z(\myexu/_2415_ ) );
BUF_X1 \myexu/_5726_ ( .A(\myexu/_0238_ ), .Z(\myexu/_2884_ ) );
BUF_X1 \myexu/_5727_ ( .A(\EX_LS_result_reg [30] ), .Z(\myexu/_2417_ ) );
BUF_X1 \myexu/_5728_ ( .A(\myexu/_0239_ ), .Z(\myexu/_2885_ ) );
BUF_X1 \myexu/_5729_ ( .A(\EX_LS_result_reg [31] ), .Z(\myexu/_2418_ ) );
BUF_X1 \myexu/_5730_ ( .A(\myexu/_0240_ ), .Z(\myexu/_2886_ ) );
BUF_X1 \myexu/_5731_ ( .A(\myexu/_0110_ ), .Z(\myexu/_2756_ ) );
BUF_X1 \myexu/_5732_ ( .A(\myexu/_0111_ ), .Z(\myexu/_2757_ ) );
BUF_X1 \myexu/_5733_ ( .A(\myexu/_0112_ ), .Z(\myexu/_2758_ ) );
BUF_X1 \myexu/_5734_ ( .A(\myexu/_0113_ ), .Z(\myexu/_2759_ ) );
BUF_X1 \myexu/_5735_ ( .A(\myexu/_0114_ ), .Z(\myexu/_2760_ ) );
BUF_X1 \myexu/_5736_ ( .A(\myexu/_0115_ ), .Z(\myexu/_2761_ ) );
BUF_X1 \myexu/_5737_ ( .A(\myexu/_0116_ ), .Z(\myexu/_2762_ ) );
BUF_X1 \myexu/_5738_ ( .A(\myexu/_0117_ ), .Z(\myexu/_2763_ ) );
BUF_X1 \myexu/_5739_ ( .A(\myexu/_0118_ ), .Z(\myexu/_2764_ ) );
BUF_X1 \myexu/_5740_ ( .A(\myexu/_0119_ ), .Z(\myexu/_2765_ ) );
BUF_X1 \myexu/_5741_ ( .A(\myexu/_0120_ ), .Z(\myexu/_2766_ ) );
BUF_X1 \myexu/_5742_ ( .A(\myexu/_0121_ ), .Z(\myexu/_2767_ ) );
BUF_X1 \myexu/_5743_ ( .A(\myexu/_0122_ ), .Z(\myexu/_2768_ ) );
BUF_X1 \myexu/_5744_ ( .A(\myexu/_0123_ ), .Z(\myexu/_2769_ ) );
BUF_X1 \myexu/_5745_ ( .A(\myexu/_0124_ ), .Z(\myexu/_2770_ ) );
BUF_X1 \myexu/_5746_ ( .A(\myexu/_0125_ ), .Z(\myexu/_2771_ ) );
BUF_X1 \myexu/_5747_ ( .A(\myexu/_0126_ ), .Z(\myexu/_2772_ ) );
BUF_X1 \myexu/_5748_ ( .A(\myexu/_0127_ ), .Z(\myexu/_2773_ ) );
BUF_X1 \myexu/_5749_ ( .A(\myexu/_0128_ ), .Z(\myexu/_2774_ ) );
BUF_X1 \myexu/_5750_ ( .A(\myexu/_0129_ ), .Z(\myexu/_2775_ ) );
BUF_X1 \myexu/_5751_ ( .A(\myexu/_0130_ ), .Z(\myexu/_2776_ ) );
BUF_X1 \myexu/_5752_ ( .A(\myexu/_0131_ ), .Z(\myexu/_2777_ ) );
BUF_X1 \myexu/_5753_ ( .A(\myexu/_0132_ ), .Z(\myexu/_2778_ ) );
BUF_X1 \myexu/_5754_ ( .A(\myexu/_0133_ ), .Z(\myexu/_2779_ ) );
BUF_X1 \myexu/_5755_ ( .A(\myexu/_0134_ ), .Z(\myexu/_2780_ ) );
BUF_X1 \myexu/_5756_ ( .A(\myexu/_0135_ ), .Z(\myexu/_2781_ ) );
BUF_X1 \myexu/_5757_ ( .A(\myexu/_0136_ ), .Z(\myexu/_2782_ ) );
BUF_X1 \myexu/_5758_ ( .A(\myexu/_0137_ ), .Z(\myexu/_2783_ ) );
BUF_X1 \myexu/_5759_ ( .A(\myexu/_0138_ ), .Z(\myexu/_2784_ ) );
BUF_X1 \myexu/_5760_ ( .A(\myexu/_0139_ ), .Z(\myexu/_2785_ ) );
BUF_X1 \myexu/_5761_ ( .A(\myexu/_0140_ ), .Z(\myexu/_2786_ ) );
BUF_X1 \myexu/_5762_ ( .A(\myexu/_0141_ ), .Z(\myexu/_2787_ ) );
BUF_X1 \myexu/_5763_ ( .A(\myexu/_0142_ ), .Z(\myexu/_2788_ ) );
BUF_X1 \myexu/_5764_ ( .A(\myexu/_0143_ ), .Z(\myexu/_2789_ ) );
BUF_X1 \myexu/_5765_ ( .A(\myexu/_0144_ ), .Z(\myexu/_2790_ ) );
BUF_X1 \myexu/_5766_ ( .A(\myexu/_0145_ ), .Z(\myexu/_2791_ ) );
BUF_X1 \myexu/_5767_ ( .A(\myexu/_0146_ ), .Z(\myexu/_2792_ ) );
BUF_X1 \myexu/_5768_ ( .A(\myexu/_0147_ ), .Z(\myexu/_2793_ ) );
BUF_X1 \myexu/_5769_ ( .A(\myexu/_0148_ ), .Z(\myexu/_2794_ ) );
BUF_X1 \myexu/_5770_ ( .A(\myexu/_0149_ ), .Z(\myexu/_2795_ ) );
BUF_X1 \myexu/_5771_ ( .A(\myexu/_0150_ ), .Z(\myexu/_2796_ ) );
BUF_X1 \myexu/_5772_ ( .A(\myexu/_0151_ ), .Z(\myexu/_2797_ ) );
BUF_X1 \myexu/_5773_ ( .A(\myexu/_0152_ ), .Z(\myexu/_2798_ ) );
BUF_X1 \myexu/_5774_ ( .A(\myexu/_0153_ ), .Z(\myexu/_2799_ ) );
BUF_X1 \myexu/_5775_ ( .A(\myexu/_0154_ ), .Z(\myexu/_2800_ ) );
BUF_X1 \myexu/_5776_ ( .A(\myexu/_0155_ ), .Z(\myexu/_2801_ ) );
BUF_X1 \myexu/_5777_ ( .A(\myexu/_0156_ ), .Z(\myexu/_2802_ ) );
BUF_X1 \myexu/_5778_ ( .A(\myexu/_0157_ ), .Z(\myexu/_2803_ ) );
BUF_X1 \myexu/_5779_ ( .A(\myexu/_0158_ ), .Z(\myexu/_2804_ ) );
BUF_X1 \myexu/_5780_ ( .A(\myexu/_0159_ ), .Z(\myexu/_2805_ ) );
BUF_X1 \myexu/_5781_ ( .A(\myexu/_0160_ ), .Z(\myexu/_2806_ ) );
BUF_X1 \myexu/_5782_ ( .A(\myexu/_0161_ ), .Z(\myexu/_2807_ ) );
BUF_X1 \myexu/_5783_ ( .A(\myexu/_0162_ ), .Z(\myexu/_2808_ ) );
BUF_X1 \myexu/_5784_ ( .A(\myexu/_0163_ ), .Z(\myexu/_2809_ ) );
BUF_X1 \myexu/_5785_ ( .A(\myexu/_0164_ ), .Z(\myexu/_2810_ ) );
BUF_X1 \myexu/_5786_ ( .A(\myexu/_0165_ ), .Z(\myexu/_2811_ ) );
BUF_X1 \myexu/_5787_ ( .A(\myexu/_0166_ ), .Z(\myexu/_2812_ ) );
BUF_X1 \myexu/_5788_ ( .A(\myexu/_0167_ ), .Z(\myexu/_2813_ ) );
BUF_X1 \myexu/_5789_ ( .A(\myexu/_0168_ ), .Z(\myexu/_2814_ ) );
BUF_X1 \myexu/_5790_ ( .A(\myexu/_0169_ ), .Z(\myexu/_2815_ ) );
BUF_X1 \myexu/_5791_ ( .A(\myexu/_0170_ ), .Z(\myexu/_2816_ ) );
BUF_X1 \myexu/_5792_ ( .A(\myexu/_0171_ ), .Z(\myexu/_2817_ ) );
BUF_X1 \myexu/_5793_ ( .A(\myexu/_0172_ ), .Z(\myexu/_2818_ ) );
BUF_X1 \myexu/_5794_ ( .A(\myexu/_0173_ ), .Z(\myexu/_2819_ ) );
BUF_X1 \myexu/_5795_ ( .A(\myexu/_0174_ ), .Z(\myexu/_2820_ ) );
BUF_X1 \myexu/_5796_ ( .A(\myexu/_0175_ ), .Z(\myexu/_2821_ ) );
BUF_X1 \myexu/_5797_ ( .A(\myexu/_0176_ ), .Z(\myexu/_2822_ ) );
BUF_X1 \myexu/_5798_ ( .A(\myexu/_0177_ ), .Z(\myexu/_2823_ ) );
BUF_X1 \myexu/_5799_ ( .A(\myexu/_0178_ ), .Z(\myexu/_2824_ ) );
BUF_X1 \myexu/_5800_ ( .A(\myexu/_0179_ ), .Z(\myexu/_2825_ ) );
BUF_X1 \myexu/_5801_ ( .A(\myexu/_0180_ ), .Z(\myexu/_2826_ ) );
BUF_X1 \myexu/_5802_ ( .A(\myexu/_0181_ ), .Z(\myexu/_2827_ ) );
BUF_X1 \myexu/_5803_ ( .A(\myexu/_0182_ ), .Z(\myexu/_2828_ ) );
BUF_X1 \myexu/_5804_ ( .A(\myexu/_0183_ ), .Z(\myexu/_2829_ ) );
BUF_X1 \myexu/_5805_ ( .A(\myexu/_0184_ ), .Z(\myexu/_2830_ ) );
BUF_X1 \myexu/_5806_ ( .A(\myexu/_0185_ ), .Z(\myexu/_2831_ ) );
BUF_X1 \myexu/_5807_ ( .A(\myexu/_0186_ ), .Z(\myexu/_2832_ ) );
BUF_X1 \myexu/_5808_ ( .A(\myexu/_0187_ ), .Z(\myexu/_2833_ ) );
BUF_X1 \myexu/_5809_ ( .A(\myexu/_0188_ ), .Z(\myexu/_2834_ ) );
AND2_X1 \myexu/myalu/_1392_ ( .A1(\myexu/myalu/_1377_ ), .A2(\myexu/myalu/_1345_ ), .ZN(\myexu/myalu/_0003_ ) );
NOR2_X1 \myexu/myalu/_1393_ ( .A1(\myexu/myalu/_1377_ ), .A2(\myexu/myalu/_1345_ ), .ZN(\myexu/myalu/_0013_ ) );
NOR2_X1 \myexu/myalu/_1394_ ( .A1(\myexu/myalu/_0003_ ), .A2(\myexu/myalu/_0013_ ), .ZN(\myexu/myalu/_0024_ ) );
XOR2_X1 \myexu/myalu/_1395_ ( .A(\myexu/myalu/_1376_ ), .B(\myexu/myalu/_1344_ ), .Z(\myexu/myalu/_0035_ ) );
XOR2_X1 \myexu/myalu/_1396_ ( .A(\myexu/myalu/_1378_ ), .B(\myexu/myalu/_1346_ ), .Z(\myexu/myalu/_0045_ ) );
AND2_X1 \myexu/myalu/_1397_ ( .A1(\myexu/myalu/_1379_ ), .A2(\myexu/myalu/_1347_ ), .ZN(\myexu/myalu/_0056_ ) );
NOR2_X1 \myexu/myalu/_1398_ ( .A1(\myexu/myalu/_1379_ ), .A2(\myexu/myalu/_1347_ ), .ZN(\myexu/myalu/_0066_ ) );
NOR2_X1 \myexu/myalu/_1399_ ( .A1(\myexu/myalu/_0056_ ), .A2(\myexu/myalu/_0066_ ), .ZN(\myexu/myalu/_0077_ ) );
OR4_X1 \myexu/myalu/_1400_ ( .A1(\myexu/myalu/_0024_ ), .A2(\myexu/myalu/_0035_ ), .A3(\myexu/myalu/_0045_ ), .A4(\myexu/myalu/_0077_ ), .ZN(\myexu/myalu/_0088_ ) );
XOR2_X1 \myexu/myalu/_1401_ ( .A(\myexu/myalu/_1384_ ), .B(\myexu/myalu/_1352_ ), .Z(\myexu/myalu/_0098_ ) );
XOR2_X1 \myexu/myalu/_1402_ ( .A(\myexu/myalu/_1383_ ), .B(\myexu/myalu/_1351_ ), .Z(\myexu/myalu/_0109_ ) );
NOR2_X1 \myexu/myalu/_1403_ ( .A1(\myexu/myalu/_0098_ ), .A2(\myexu/myalu/_0109_ ), .ZN(\myexu/myalu/_0119_ ) );
AND2_X1 \myexu/myalu/_1404_ ( .A1(\myexu/myalu/_1381_ ), .A2(\myexu/myalu/_1349_ ), .ZN(\myexu/myalu/_0130_ ) );
NOR2_X1 \myexu/myalu/_1405_ ( .A1(\myexu/myalu/_1381_ ), .A2(\myexu/myalu/_1349_ ), .ZN(\myexu/myalu/_0141_ ) );
NOR2_X1 \myexu/myalu/_1406_ ( .A1(\myexu/myalu/_0130_ ), .A2(\myexu/myalu/_0141_ ), .ZN(\myexu/myalu/_0152_ ) );
INV_X1 \myexu/myalu/_1407_ ( .A(\myexu/myalu/_0152_ ), .ZN(\myexu/myalu/_0162_ ) );
XOR2_X1 \myexu/myalu/_1408_ ( .A(\myexu/myalu/_1380_ ), .B(\myexu/myalu/_1348_ ), .Z(\myexu/myalu/_0173_ ) );
INV_X1 \myexu/myalu/_1409_ ( .A(\myexu/myalu/_0173_ ), .ZN(\myexu/myalu/_0183_ ) );
NAND3_X1 \myexu/myalu/_1410_ ( .A1(\myexu/myalu/_0119_ ), .A2(\myexu/myalu/_0162_ ), .A3(\myexu/myalu/_0183_ ), .ZN(\myexu/myalu/_0194_ ) );
NOR2_X1 \myexu/myalu/_1411_ ( .A1(\myexu/myalu/_0088_ ), .A2(\myexu/myalu/_0194_ ), .ZN(\myexu/myalu/_0204_ ) );
XOR2_X1 \myexu/myalu/_1412_ ( .A(\myexu/myalu/_1374_ ), .B(\myexu/myalu/_1342_ ), .Z(\myexu/myalu/_0215_ ) );
AND2_X1 \myexu/myalu/_1413_ ( .A1(\myexu/myalu/_1375_ ), .A2(\myexu/myalu/_1343_ ), .ZN(\myexu/myalu/_0226_ ) );
NOR2_X1 \myexu/myalu/_1414_ ( .A1(\myexu/myalu/_1375_ ), .A2(\myexu/myalu/_1343_ ), .ZN(\myexu/myalu/_0236_ ) );
NOR2_X1 \myexu/myalu/_1415_ ( .A1(\myexu/myalu/_0226_ ), .A2(\myexu/myalu/_0236_ ), .ZN(\myexu/myalu/_0247_ ) );
NOR2_X1 \myexu/myalu/_1416_ ( .A1(\myexu/myalu/_0215_ ), .A2(\myexu/myalu/_0247_ ), .ZN(\myexu/myalu/_0258_ ) );
XOR2_X1 \myexu/myalu/_1417_ ( .A(\myexu/myalu/_1372_ ), .B(\myexu/myalu/_1340_ ), .Z(\myexu/myalu/_0268_ ) );
AND2_X1 \myexu/myalu/_1418_ ( .A1(\myexu/myalu/_1373_ ), .A2(\myexu/myalu/_1341_ ), .ZN(\myexu/myalu/_0279_ ) );
NOR2_X1 \myexu/myalu/_1419_ ( .A1(\myexu/myalu/_1373_ ), .A2(\myexu/myalu/_1341_ ), .ZN(\myexu/myalu/_0290_ ) );
NOR2_X1 \myexu/myalu/_1420_ ( .A1(\myexu/myalu/_0279_ ), .A2(\myexu/myalu/_0290_ ), .ZN(\myexu/myalu/_0301_ ) );
NOR2_X1 \myexu/myalu/_1421_ ( .A1(\myexu/myalu/_0268_ ), .A2(\myexu/myalu/_0301_ ), .ZN(\myexu/myalu/_0311_ ) );
XOR2_X1 \myexu/myalu/_1422_ ( .A(\myexu/myalu/_1369_ ), .B(\myexu/myalu/_1337_ ), .Z(\myexu/myalu/_0322_ ) );
AND2_X1 \myexu/myalu/_1423_ ( .A1(\myexu/myalu/_1370_ ), .A2(\myexu/myalu/_1338_ ), .ZN(\myexu/myalu/_0333_ ) );
NOR2_X1 \myexu/myalu/_1424_ ( .A1(\myexu/myalu/_1370_ ), .A2(\myexu/myalu/_1338_ ), .ZN(\myexu/myalu/_0343_ ) );
NOR2_X1 \myexu/myalu/_1425_ ( .A1(\myexu/myalu/_0333_ ), .A2(\myexu/myalu/_0343_ ), .ZN(\myexu/myalu/_0354_ ) );
NOR2_X1 \myexu/myalu/_1426_ ( .A1(\myexu/myalu/_0322_ ), .A2(\myexu/myalu/_0354_ ), .ZN(\myexu/myalu/_0364_ ) );
NAND3_X1 \myexu/myalu/_1427_ ( .A1(\myexu/myalu/_0258_ ), .A2(\myexu/myalu/_0311_ ), .A3(\myexu/myalu/_0364_ ), .ZN(\myexu/myalu/_0375_ ) );
AND2_X2 \myexu/myalu/_1428_ ( .A1(\myexu/myalu/_1368_ ), .A2(\myexu/myalu/_1336_ ), .ZN(\myexu/myalu/_0385_ ) );
NOR2_X1 \myexu/myalu/_1429_ ( .A1(\myexu/myalu/_1368_ ), .A2(\myexu/myalu/_1336_ ), .ZN(\myexu/myalu/_0396_ ) );
NOR2_X1 \myexu/myalu/_1430_ ( .A1(\myexu/myalu/_0385_ ), .A2(\myexu/myalu/_0396_ ), .ZN(\myexu/myalu/_0407_ ) );
XOR2_X1 \myexu/myalu/_1431_ ( .A(\myexu/myalu/_1367_ ), .B(\myexu/myalu/_1335_ ), .Z(\myexu/myalu/_0417_ ) );
OR3_X1 \myexu/myalu/_1432_ ( .A1(\myexu/myalu/_0375_ ), .A2(\myexu/myalu/_0407_ ), .A3(\myexu/myalu/_0417_ ), .ZN(\myexu/myalu/_0428_ ) );
XOR2_X1 \myexu/myalu/_1433_ ( .A(\myexu/myalu/_1365_ ), .B(\myexu/myalu/_1333_ ), .Z(\myexu/myalu/_0438_ ) );
AND2_X4 \myexu/myalu/_1434_ ( .A1(\myexu/myalu/_1366_ ), .A2(\myexu/myalu/_1334_ ), .ZN(\myexu/myalu/_0449_ ) );
NOR2_X1 \myexu/myalu/_1435_ ( .A1(\myexu/myalu/_1366_ ), .A2(\myexu/myalu/_1334_ ), .ZN(\myexu/myalu/_0454_ ) );
NOR2_X1 \myexu/myalu/_1436_ ( .A1(\myexu/myalu/_0449_ ), .A2(\myexu/myalu/_0454_ ), .ZN(\myexu/myalu/_0455_ ) );
NOR2_X1 \myexu/myalu/_1437_ ( .A1(\myexu/myalu/_0438_ ), .A2(\myexu/myalu/_0455_ ), .ZN(\myexu/myalu/_0456_ ) );
AND2_X1 \myexu/myalu/_1438_ ( .A1(\myexu/myalu/_1364_ ), .A2(\myexu/myalu/_1332_ ), .ZN(\myexu/myalu/_0457_ ) );
NOR2_X1 \myexu/myalu/_1439_ ( .A1(\myexu/myalu/_1364_ ), .A2(\myexu/myalu/_1332_ ), .ZN(\myexu/myalu/_0458_ ) );
NOR2_X2 \myexu/myalu/_1440_ ( .A1(\myexu/myalu/_0457_ ), .A2(\myexu/myalu/_0458_ ), .ZN(\myexu/myalu/_0459_ ) );
INV_X1 \myexu/myalu/_1441_ ( .A(\myexu/myalu/_0459_ ), .ZN(\myexu/myalu/_0460_ ) );
XOR2_X1 \myexu/myalu/_1442_ ( .A(\myexu/myalu/_1363_ ), .B(\myexu/myalu/_1331_ ), .Z(\myexu/myalu/_0461_ ) );
INV_X1 \myexu/myalu/_1443_ ( .A(\myexu/myalu/_0461_ ), .ZN(\myexu/myalu/_0462_ ) );
AND3_X1 \myexu/myalu/_1444_ ( .A1(\myexu/myalu/_0456_ ), .A2(\myexu/myalu/_0460_ ), .A3(\myexu/myalu/_0462_ ), .ZN(\myexu/myalu/_0463_ ) );
XOR2_X2 \myexu/myalu/_1445_ ( .A(\myexu/myalu/_1361_ ), .B(\myexu/myalu/_1329_ ), .Z(\myexu/myalu/_0464_ ) );
AND2_X1 \myexu/myalu/_1446_ ( .A1(\myexu/myalu/_1362_ ), .A2(\myexu/myalu/_1330_ ), .ZN(\myexu/myalu/_0465_ ) );
NOR2_X2 \myexu/myalu/_1447_ ( .A1(\myexu/myalu/_1362_ ), .A2(\myexu/myalu/_1330_ ), .ZN(\myexu/myalu/_0466_ ) );
NOR2_X1 \myexu/myalu/_1448_ ( .A1(\myexu/myalu/_0465_ ), .A2(\myexu/myalu/_0466_ ), .ZN(\myexu/myalu/_0467_ ) );
NOR2_X1 \myexu/myalu/_1449_ ( .A1(\myexu/myalu/_0464_ ), .A2(\myexu/myalu/_0467_ ), .ZN(\myexu/myalu/_0468_ ) );
AND2_X1 \myexu/myalu/_1450_ ( .A1(\myexu/myalu/_1391_ ), .A2(\myexu/myalu/_1359_ ), .ZN(\myexu/myalu/_0469_ ) );
NOR2_X1 \myexu/myalu/_1451_ ( .A1(\myexu/myalu/_1391_ ), .A2(\myexu/myalu/_1359_ ), .ZN(\myexu/myalu/_0470_ ) );
NOR2_X1 \myexu/myalu/_1452_ ( .A1(\myexu/myalu/_0469_ ), .A2(\myexu/myalu/_0470_ ), .ZN(\myexu/myalu/_0471_ ) );
INV_X1 \myexu/myalu/_1453_ ( .A(\myexu/myalu/_0471_ ), .ZN(\myexu/myalu/_0472_ ) );
XOR2_X1 \myexu/myalu/_1454_ ( .A(\myexu/myalu/_1390_ ), .B(\myexu/myalu/_1358_ ), .Z(\myexu/myalu/_0473_ ) );
INV_X1 \myexu/myalu/_1455_ ( .A(\myexu/myalu/_0473_ ), .ZN(\myexu/myalu/_0474_ ) );
AND4_X1 \myexu/myalu/_1456_ ( .A1(\myexu/myalu/_0463_ ), .A2(\myexu/myalu/_0468_ ), .A3(\myexu/myalu/_0472_ ), .A4(\myexu/myalu/_0474_ ), .ZN(\myexu/myalu/_0475_ ) );
INV_X1 \myexu/myalu/_1457_ ( .A(\myexu/myalu/_1356_ ), .ZN(\myexu/myalu/_0476_ ) );
NOR2_X1 \myexu/myalu/_1458_ ( .A1(\myexu/myalu/_0476_ ), .A2(\myexu/myalu/_1388_ ), .ZN(\myexu/myalu/_0477_ ) );
AND2_X4 \myexu/myalu/_1459_ ( .A1(\myexu/myalu/_1389_ ), .A2(\myexu/myalu/_1357_ ), .ZN(\myexu/myalu/_0478_ ) );
NOR2_X1 \myexu/myalu/_1460_ ( .A1(\myexu/myalu/_1389_ ), .A2(\myexu/myalu/_1357_ ), .ZN(\myexu/myalu/_0479_ ) );
OAI21_X1 \myexu/myalu/_1461_ ( .A(\myexu/myalu/_0477_ ), .B1(\myexu/myalu/_0478_ ), .B2(\myexu/myalu/_0479_ ), .ZN(\myexu/myalu/_0480_ ) );
INV_X1 \myexu/myalu/_1462_ ( .A(\myexu/myalu/_1357_ ), .ZN(\myexu/myalu/_0481_ ) );
XOR2_X2 \myexu/myalu/_1463_ ( .A(\myexu/myalu/_1387_ ), .B(\myexu/myalu/_1355_ ), .Z(\myexu/myalu/_0482_ ) );
INV_X1 \myexu/myalu/_1464_ ( .A(\myexu/myalu/_1354_ ), .ZN(\myexu/myalu/_0483_ ) );
NOR3_X1 \myexu/myalu/_1465_ ( .A1(\myexu/myalu/_0482_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0483_ ), .ZN(\myexu/myalu/_0484_ ) );
INV_X1 \myexu/myalu/_1466_ ( .A(\myexu/myalu/_1387_ ), .ZN(\myexu/myalu/_0485_ ) );
AOI21_X1 \myexu/myalu/_1467_ ( .A(\myexu/myalu/_0484_ ), .B1(\myexu/myalu/_0485_ ), .B2(\myexu/myalu/_1355_ ), .ZN(\myexu/myalu/_0486_ ) );
XOR2_X1 \myexu/myalu/_1468_ ( .A(\myexu/myalu/_1388_ ), .B(\myexu/myalu/_1356_ ), .Z(\myexu/myalu/_0487_ ) );
NOR2_X2 \myexu/myalu/_1469_ ( .A1(\myexu/myalu/_0478_ ), .A2(\myexu/myalu/_0479_ ), .ZN(\myexu/myalu/_0488_ ) );
OR2_X1 \myexu/myalu/_1470_ ( .A1(\myexu/myalu/_0487_ ), .A2(\myexu/myalu/_0488_ ), .ZN(\myexu/myalu/_0489_ ) );
OAI221_X1 \myexu/myalu/_1471_ ( .A(\myexu/myalu/_0480_ ), .B1(\myexu/myalu/_1389_ ), .B2(\myexu/myalu/_0481_ ), .C1(\myexu/myalu/_0486_ ), .C2(\myexu/myalu/_0489_ ), .ZN(\myexu/myalu/_0490_ ) );
XOR2_X1 \myexu/myalu/_1472_ ( .A(fanout_net_17 ), .B(\myexu/myalu/_1354_ ), .Z(\myexu/myalu/_0491_ ) );
OR4_X1 \myexu/myalu/_1473_ ( .A1(\myexu/myalu/_0488_ ), .A2(\myexu/myalu/_0487_ ), .A3(\myexu/myalu/_0482_ ), .A4(\myexu/myalu/_0491_ ), .ZN(\myexu/myalu/_0492_ ) );
XNOR2_X1 \myexu/myalu/_1474_ ( .A(fanout_net_15 ), .B(\myexu/myalu/_1353_ ), .ZN(\myexu/myalu/_0493_ ) );
XOR2_X1 \myexu/myalu/_1475_ ( .A(fanout_net_13 ), .B(\myexu/myalu/_1350_ ), .Z(\myexu/myalu/_0494_ ) );
INV_X1 \myexu/myalu/_1476_ ( .A(\myexu/myalu/_0494_ ), .ZN(\myexu/myalu/_0495_ ) );
XOR2_X2 \myexu/myalu/_1477_ ( .A(fanout_net_11 ), .B(\myexu/myalu/_1339_ ), .Z(\myexu/myalu/_0496_ ) );
INV_X1 \myexu/myalu/_1478_ ( .A(\myexu/myalu/_1328_ ), .ZN(\myexu/myalu/_0497_ ) );
AOI21_X1 \myexu/myalu/_1479_ ( .A(\myexu/myalu/_0496_ ), .B1(fanout_net_9 ), .B2(\myexu/myalu/_0497_ ), .ZN(\myexu/myalu/_0498_ ) );
INV_X1 \myexu/myalu/_1480_ ( .A(\myexu/myalu/_1339_ ), .ZN(\myexu/myalu/_0499_ ) );
NOR2_X1 \myexu/myalu/_1481_ ( .A1(\myexu/myalu/_0499_ ), .A2(fanout_net_11 ), .ZN(\myexu/myalu/_0500_ ) );
OAI211_X2 \myexu/myalu/_1482_ ( .A(\myexu/myalu/_0493_ ), .B(\myexu/myalu/_0495_ ), .C1(\myexu/myalu/_0498_ ), .C2(\myexu/myalu/_0500_ ), .ZN(\myexu/myalu/_0501_ ) );
INV_X1 \myexu/myalu/_1483_ ( .A(\myexu/myalu/_1350_ ), .ZN(\myexu/myalu/_0502_ ) );
NOR2_X1 \myexu/myalu/_1484_ ( .A1(\myexu/myalu/_0502_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0503_ ) );
AND2_X1 \myexu/myalu/_1485_ ( .A1(\myexu/myalu/_0493_ ), .A2(\myexu/myalu/_0503_ ), .ZN(\myexu/myalu/_0504_ ) );
INV_X32 \myexu/myalu/_1486_ ( .A(fanout_net_15 ), .ZN(\myexu/myalu/_0505_ ) );
BUF_X4 \myexu/myalu/_1487_ ( .A(\myexu/myalu/_0505_ ), .Z(\myexu/myalu/_0506_ ) );
AOI21_X1 \myexu/myalu/_1488_ ( .A(\myexu/myalu/_0504_ ), .B1(\myexu/myalu/_0506_ ), .B2(\myexu/myalu/_1353_ ), .ZN(\myexu/myalu/_0507_ ) );
AOI21_X1 \myexu/myalu/_1489_ ( .A(\myexu/myalu/_0492_ ), .B1(\myexu/myalu/_0501_ ), .B2(\myexu/myalu/_0507_ ), .ZN(\myexu/myalu/_0508_ ) );
OAI21_X1 \myexu/myalu/_1490_ ( .A(\myexu/myalu/_0475_ ), .B1(\myexu/myalu/_0490_ ), .B2(\myexu/myalu/_0508_ ), .ZN(\myexu/myalu/_0509_ ) );
INV_X1 \myexu/myalu/_1491_ ( .A(\myexu/myalu/_1358_ ), .ZN(\myexu/myalu/_0510_ ) );
NOR3_X1 \myexu/myalu/_1492_ ( .A1(\myexu/myalu/_0471_ ), .A2(\myexu/myalu/_1390_ ), .A3(\myexu/myalu/_0510_ ), .ZN(\myexu/myalu/_0511_ ) );
INV_X1 \myexu/myalu/_1493_ ( .A(\myexu/myalu/_1359_ ), .ZN(\myexu/myalu/_0512_ ) );
NOR2_X1 \myexu/myalu/_1494_ ( .A1(\myexu/myalu/_0512_ ), .A2(\myexu/myalu/_1391_ ), .ZN(\myexu/myalu/_0513_ ) );
OAI21_X1 \myexu/myalu/_1495_ ( .A(\myexu/myalu/_0468_ ), .B1(\myexu/myalu/_0511_ ), .B2(\myexu/myalu/_0513_ ), .ZN(\myexu/myalu/_0514_ ) );
INV_X1 \myexu/myalu/_1496_ ( .A(\myexu/myalu/_1329_ ), .ZN(\myexu/myalu/_0515_ ) );
OR3_X1 \myexu/myalu/_1497_ ( .A1(\myexu/myalu/_0467_ ), .A2(\myexu/myalu/_1361_ ), .A3(\myexu/myalu/_0515_ ), .ZN(\myexu/myalu/_0516_ ) );
INV_X1 \myexu/myalu/_1498_ ( .A(\myexu/myalu/_1362_ ), .ZN(\myexu/myalu/_0517_ ) );
NAND2_X1 \myexu/myalu/_1499_ ( .A1(\myexu/myalu/_0517_ ), .A2(\myexu/myalu/_1330_ ), .ZN(\myexu/myalu/_0518_ ) );
NAND3_X1 \myexu/myalu/_1500_ ( .A1(\myexu/myalu/_0514_ ), .A2(\myexu/myalu/_0516_ ), .A3(\myexu/myalu/_0518_ ), .ZN(\myexu/myalu/_0519_ ) );
NAND2_X1 \myexu/myalu/_1501_ ( .A1(\myexu/myalu/_0519_ ), .A2(\myexu/myalu/_0463_ ), .ZN(\myexu/myalu/_0520_ ) );
INV_X1 \myexu/myalu/_1502_ ( .A(\myexu/myalu/_1331_ ), .ZN(\myexu/myalu/_0521_ ) );
NOR3_X1 \myexu/myalu/_1503_ ( .A1(\myexu/myalu/_0459_ ), .A2(\myexu/myalu/_1363_ ), .A3(\myexu/myalu/_0521_ ), .ZN(\myexu/myalu/_0522_ ) );
INV_X1 \myexu/myalu/_1504_ ( .A(\myexu/myalu/_1332_ ), .ZN(\myexu/myalu/_0523_ ) );
NOR2_X1 \myexu/myalu/_1505_ ( .A1(\myexu/myalu/_0523_ ), .A2(\myexu/myalu/_1364_ ), .ZN(\myexu/myalu/_0524_ ) );
OAI21_X1 \myexu/myalu/_1506_ ( .A(\myexu/myalu/_0456_ ), .B1(\myexu/myalu/_0522_ ), .B2(\myexu/myalu/_0524_ ), .ZN(\myexu/myalu/_0525_ ) );
INV_X1 \myexu/myalu/_1507_ ( .A(\myexu/myalu/_1333_ ), .ZN(\myexu/myalu/_0526_ ) );
OR3_X1 \myexu/myalu/_1508_ ( .A1(\myexu/myalu/_0455_ ), .A2(\myexu/myalu/_1365_ ), .A3(\myexu/myalu/_0526_ ), .ZN(\myexu/myalu/_0527_ ) );
INV_X1 \myexu/myalu/_1509_ ( .A(\myexu/myalu/_1366_ ), .ZN(\myexu/myalu/_0528_ ) );
NAND2_X1 \myexu/myalu/_1510_ ( .A1(\myexu/myalu/_0528_ ), .A2(\myexu/myalu/_1334_ ), .ZN(\myexu/myalu/_0529_ ) );
AND3_X1 \myexu/myalu/_1511_ ( .A1(\myexu/myalu/_0525_ ), .A2(\myexu/myalu/_0527_ ), .A3(\myexu/myalu/_0529_ ), .ZN(\myexu/myalu/_0530_ ) );
AND2_X1 \myexu/myalu/_1512_ ( .A1(\myexu/myalu/_0520_ ), .A2(\myexu/myalu/_0530_ ), .ZN(\myexu/myalu/_0531_ ) );
AOI21_X1 \myexu/myalu/_1513_ ( .A(\myexu/myalu/_0428_ ), .B1(\myexu/myalu/_0509_ ), .B2(\myexu/myalu/_0531_ ), .ZN(\myexu/myalu/_0532_ ) );
AND2_X1 \myexu/myalu/_1514_ ( .A1(\myexu/myalu/_0258_ ), .A2(\myexu/myalu/_0311_ ), .ZN(\myexu/myalu/_0533_ ) );
INV_X1 \myexu/myalu/_1515_ ( .A(\myexu/myalu/_1335_ ), .ZN(\myexu/myalu/_0534_ ) );
NOR3_X1 \myexu/myalu/_1516_ ( .A1(\myexu/myalu/_0407_ ), .A2(\myexu/myalu/_1367_ ), .A3(\myexu/myalu/_0534_ ), .ZN(\myexu/myalu/_0535_ ) );
INV_X1 \myexu/myalu/_1517_ ( .A(\myexu/myalu/_1336_ ), .ZN(\myexu/myalu/_0536_ ) );
NOR2_X1 \myexu/myalu/_1518_ ( .A1(\myexu/myalu/_0536_ ), .A2(\myexu/myalu/_1368_ ), .ZN(\myexu/myalu/_0537_ ) );
OAI21_X1 \myexu/myalu/_1519_ ( .A(\myexu/myalu/_0364_ ), .B1(\myexu/myalu/_0535_ ), .B2(\myexu/myalu/_0537_ ), .ZN(\myexu/myalu/_0538_ ) );
INV_X1 \myexu/myalu/_1520_ ( .A(\myexu/myalu/_1370_ ), .ZN(\myexu/myalu/_0539_ ) );
NAND2_X1 \myexu/myalu/_1521_ ( .A1(\myexu/myalu/_0539_ ), .A2(\myexu/myalu/_1338_ ), .ZN(\myexu/myalu/_0540_ ) );
NAND2_X1 \myexu/myalu/_1522_ ( .A1(\myexu/myalu/_0538_ ), .A2(\myexu/myalu/_0540_ ), .ZN(\myexu/myalu/_0541_ ) );
INV_X1 \myexu/myalu/_1523_ ( .A(\myexu/myalu/_1337_ ), .ZN(\myexu/myalu/_0542_ ) );
NOR3_X1 \myexu/myalu/_1524_ ( .A1(\myexu/myalu/_0354_ ), .A2(\myexu/myalu/_1369_ ), .A3(\myexu/myalu/_0542_ ), .ZN(\myexu/myalu/_0543_ ) );
OAI21_X1 \myexu/myalu/_1525_ ( .A(\myexu/myalu/_0533_ ), .B1(\myexu/myalu/_0541_ ), .B2(\myexu/myalu/_0543_ ), .ZN(\myexu/myalu/_0544_ ) );
INV_X1 \myexu/myalu/_1526_ ( .A(\myexu/myalu/_1342_ ), .ZN(\myexu/myalu/_0545_ ) );
NOR3_X1 \myexu/myalu/_1527_ ( .A1(\myexu/myalu/_0247_ ), .A2(\myexu/myalu/_1374_ ), .A3(\myexu/myalu/_0545_ ), .ZN(\myexu/myalu/_0546_ ) );
INV_X1 \myexu/myalu/_1528_ ( .A(\myexu/myalu/_1375_ ), .ZN(\myexu/myalu/_0547_ ) );
AOI21_X1 \myexu/myalu/_1529_ ( .A(\myexu/myalu/_0546_ ), .B1(\myexu/myalu/_0547_ ), .B2(\myexu/myalu/_1343_ ), .ZN(\myexu/myalu/_0548_ ) );
INV_X1 \myexu/myalu/_1530_ ( .A(\myexu/myalu/_1340_ ), .ZN(\myexu/myalu/_0549_ ) );
NOR3_X1 \myexu/myalu/_1531_ ( .A1(\myexu/myalu/_0301_ ), .A2(\myexu/myalu/_1372_ ), .A3(\myexu/myalu/_0549_ ), .ZN(\myexu/myalu/_0550_ ) );
INV_X1 \myexu/myalu/_1532_ ( .A(\myexu/myalu/_1341_ ), .ZN(\myexu/myalu/_0551_ ) );
NOR2_X1 \myexu/myalu/_1533_ ( .A1(\myexu/myalu/_0551_ ), .A2(\myexu/myalu/_1373_ ), .ZN(\myexu/myalu/_0552_ ) );
OAI21_X1 \myexu/myalu/_1534_ ( .A(\myexu/myalu/_0258_ ), .B1(\myexu/myalu/_0550_ ), .B2(\myexu/myalu/_0552_ ), .ZN(\myexu/myalu/_0553_ ) );
NAND3_X1 \myexu/myalu/_1535_ ( .A1(\myexu/myalu/_0544_ ), .A2(\myexu/myalu/_0548_ ), .A3(\myexu/myalu/_0553_ ), .ZN(\myexu/myalu/_0554_ ) );
OAI21_X1 \myexu/myalu/_1536_ ( .A(\myexu/myalu/_0204_ ), .B1(\myexu/myalu/_0532_ ), .B2(\myexu/myalu/_0554_ ), .ZN(\myexu/myalu/_0555_ ) );
INV_X1 \myexu/myalu/_1537_ ( .A(\myexu/myalu/_0098_ ), .ZN(\myexu/myalu/_0556_ ) );
INV_X1 \myexu/myalu/_1538_ ( .A(\myexu/myalu/_1383_ ), .ZN(\myexu/myalu/_0557_ ) );
NAND3_X1 \myexu/myalu/_1539_ ( .A1(\myexu/myalu/_0556_ ), .A2(\myexu/myalu/_0557_ ), .A3(\myexu/myalu/_1351_ ), .ZN(\myexu/myalu/_0558_ ) );
NOR2_X1 \myexu/myalu/_1540_ ( .A1(\myexu/myalu/_0001_ ), .A2(\myexu/myalu/_0000_ ), .ZN(\myexu/myalu/_0559_ ) );
OR2_X1 \myexu/myalu/_1541_ ( .A1(\myexu/myalu/_0045_ ), .A2(\myexu/myalu/_0077_ ), .ZN(\myexu/myalu/_0560_ ) );
INV_X1 \myexu/myalu/_1542_ ( .A(\myexu/myalu/_1376_ ), .ZN(\myexu/myalu/_0561_ ) );
OAI211_X2 \myexu/myalu/_1543_ ( .A(\myexu/myalu/_0561_ ), .B(\myexu/myalu/_1344_ ), .C1(\myexu/myalu/_0003_ ), .C2(\myexu/myalu/_0013_ ), .ZN(\myexu/myalu/_0562_ ) );
INV_X1 \myexu/myalu/_1544_ ( .A(\myexu/myalu/_1377_ ), .ZN(\myexu/myalu/_0563_ ) );
NAND2_X1 \myexu/myalu/_1545_ ( .A1(\myexu/myalu/_0563_ ), .A2(\myexu/myalu/_1345_ ), .ZN(\myexu/myalu/_0564_ ) );
AOI21_X1 \myexu/myalu/_1546_ ( .A(\myexu/myalu/_0560_ ), .B1(\myexu/myalu/_0562_ ), .B2(\myexu/myalu/_0564_ ), .ZN(\myexu/myalu/_0565_ ) );
INV_X1 \myexu/myalu/_1547_ ( .A(\myexu/myalu/_1346_ ), .ZN(\myexu/myalu/_0566_ ) );
NOR3_X1 \myexu/myalu/_1548_ ( .A1(\myexu/myalu/_0077_ ), .A2(\myexu/myalu/_1378_ ), .A3(\myexu/myalu/_0566_ ), .ZN(\myexu/myalu/_0567_ ) );
INV_X1 \myexu/myalu/_1549_ ( .A(\myexu/myalu/_1347_ ), .ZN(\myexu/myalu/_0568_ ) );
NOR2_X1 \myexu/myalu/_1550_ ( .A1(\myexu/myalu/_0568_ ), .A2(\myexu/myalu/_1379_ ), .ZN(\myexu/myalu/_0569_ ) );
NOR3_X1 \myexu/myalu/_1551_ ( .A1(\myexu/myalu/_0565_ ), .A2(\myexu/myalu/_0567_ ), .A3(\myexu/myalu/_0569_ ), .ZN(\myexu/myalu/_0570_ ) );
OR2_X1 \myexu/myalu/_1552_ ( .A1(\myexu/myalu/_0570_ ), .A2(\myexu/myalu/_0194_ ), .ZN(\myexu/myalu/_0571_ ) );
INV_X1 \myexu/myalu/_1553_ ( .A(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0572_ ) );
INV_X1 \myexu/myalu/_1554_ ( .A(\myexu/myalu/_1384_ ), .ZN(\myexu/myalu/_0573_ ) );
AOI21_X1 \myexu/myalu/_1555_ ( .A(\myexu/myalu/_0572_ ), .B1(\myexu/myalu/_0573_ ), .B2(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_0574_ ) );
INV_X1 \myexu/myalu/_1556_ ( .A(\myexu/myalu/_1348_ ), .ZN(\myexu/myalu/_0575_ ) );
NOR3_X1 \myexu/myalu/_1557_ ( .A1(\myexu/myalu/_0152_ ), .A2(\myexu/myalu/_1380_ ), .A3(\myexu/myalu/_0575_ ), .ZN(\myexu/myalu/_0576_ ) );
INV_X1 \myexu/myalu/_1558_ ( .A(\myexu/myalu/_1349_ ), .ZN(\myexu/myalu/_0577_ ) );
NOR2_X1 \myexu/myalu/_1559_ ( .A1(\myexu/myalu/_0577_ ), .A2(\myexu/myalu/_1381_ ), .ZN(\myexu/myalu/_0578_ ) );
OAI21_X1 \myexu/myalu/_1560_ ( .A(\myexu/myalu/_0119_ ), .B1(\myexu/myalu/_0576_ ), .B2(\myexu/myalu/_0578_ ), .ZN(\myexu/myalu/_0579_ ) );
AND4_X1 \myexu/myalu/_1561_ ( .A1(\myexu/myalu/_0559_ ), .A2(\myexu/myalu/_0571_ ), .A3(\myexu/myalu/_0574_ ), .A4(\myexu/myalu/_0579_ ), .ZN(\myexu/myalu/_0580_ ) );
AND3_X1 \myexu/myalu/_1562_ ( .A1(\myexu/myalu/_0555_ ), .A2(\myexu/myalu/_0558_ ), .A3(\myexu/myalu/_0580_ ), .ZN(\myexu/myalu/_0581_ ) );
AND2_X1 \myexu/myalu/_1563_ ( .A1(\myexu/myalu/_1390_ ), .A2(\myexu/myalu/_1391_ ), .ZN(\myexu/myalu/_0582_ ) );
NOR2_X1 \myexu/myalu/_1564_ ( .A1(\myexu/myalu/_1390_ ), .A2(\myexu/myalu/_1391_ ), .ZN(\myexu/myalu/_0583_ ) );
NOR2_X4 \myexu/myalu/_1565_ ( .A1(fanout_net_9 ), .A2(fanout_net_11 ), .ZN(\myexu/myalu/_0584_ ) );
INV_X32 \myexu/myalu/_1566_ ( .A(fanout_net_13 ), .ZN(\myexu/myalu/_0585_ ) );
AND2_X4 \myexu/myalu/_1567_ ( .A1(\myexu/myalu/_0584_ ), .A2(\myexu/myalu/_0585_ ), .ZN(\myexu/myalu/_0586_ ) );
AND2_X4 \myexu/myalu/_1568_ ( .A1(\myexu/myalu/_0586_ ), .A2(\myexu/myalu/_0505_ ), .ZN(\myexu/myalu/_0587_ ) );
INV_X1 \myexu/myalu/_1569_ ( .A(fanout_net_17 ), .ZN(\myexu/myalu/_0588_ ) );
AND2_X4 \myexu/myalu/_1570_ ( .A1(\myexu/myalu/_0587_ ), .A2(\myexu/myalu/_0588_ ), .ZN(\myexu/myalu/_0589_ ) );
INV_X4 \myexu/myalu/_1571_ ( .A(\myexu/myalu/_0589_ ), .ZN(\myexu/myalu/_0590_ ) );
AOI21_X4 \myexu/myalu/_1572_ ( .A(\myexu/myalu/_1388_ ), .B1(\myexu/myalu/_0590_ ), .B2(\myexu/myalu/_1387_ ), .ZN(\myexu/myalu/_0591_ ) );
INV_X1 \myexu/myalu/_1573_ ( .A(\myexu/myalu/_1389_ ), .ZN(\myexu/myalu/_0592_ ) );
AND2_X4 \myexu/myalu/_1574_ ( .A1(\myexu/myalu/_0591_ ), .A2(\myexu/myalu/_0592_ ), .ZN(\myexu/myalu/_0593_ ) );
MUX2_X1 \myexu/myalu/_1575_ ( .A(\myexu/myalu/_0582_ ), .B(\myexu/myalu/_0583_ ), .S(\myexu/myalu/_0593_ ), .Z(\myexu/myalu/_0594_ ) );
NAND4_X1 \myexu/myalu/_1576_ ( .A1(\myexu/myalu/_0590_ ), .A2(\myexu/myalu/_1387_ ), .A3(\myexu/myalu/_1388_ ), .A4(\myexu/myalu/_1389_ ), .ZN(\myexu/myalu/_0595_ ) );
INV_X1 \myexu/myalu/_1577_ ( .A(\myexu/myalu/_0595_ ), .ZN(\myexu/myalu/_0596_ ) );
OAI211_X2 \myexu/myalu/_1578_ ( .A(\myexu/myalu/_0594_ ), .B(\myexu/myalu/_1352_ ), .C1(\myexu/myalu/_0593_ ), .C2(\myexu/myalu/_0596_ ), .ZN(\myexu/myalu/_0597_ ) );
AND2_X4 \myexu/myalu/_1579_ ( .A1(\myexu/myalu/_0593_ ), .A2(\myexu/myalu/_0583_ ), .ZN(\myexu/myalu/_0598_ ) );
NOR2_X1 \myexu/myalu/_1580_ ( .A1(\myexu/myalu/_1361_ ), .A2(\myexu/myalu/_1362_ ), .ZN(\myexu/myalu/_0599_ ) );
AND2_X4 \myexu/myalu/_1581_ ( .A1(\myexu/myalu/_0598_ ), .A2(\myexu/myalu/_0599_ ), .ZN(\myexu/myalu/_0600_ ) );
INV_X4 \myexu/myalu/_1582_ ( .A(\myexu/myalu/_0600_ ), .ZN(\myexu/myalu/_0601_ ) );
INV_X1 \myexu/myalu/_1583_ ( .A(\myexu/myalu/_0598_ ), .ZN(\myexu/myalu/_0602_ ) );
AND2_X1 \myexu/myalu/_1584_ ( .A1(\myexu/myalu/_1361_ ), .A2(\myexu/myalu/_1362_ ), .ZN(\myexu/myalu/_0603_ ) );
NAND2_X1 \myexu/myalu/_1585_ ( .A1(\myexu/myalu/_0602_ ), .A2(\myexu/myalu/_0603_ ), .ZN(\myexu/myalu/_0604_ ) );
AOI21_X1 \myexu/myalu/_1586_ ( .A(\myexu/myalu/_0597_ ), .B1(\myexu/myalu/_0601_ ), .B2(\myexu/myalu/_0604_ ), .ZN(\myexu/myalu/_0605_ ) );
NOR2_X4 \myexu/myalu/_1587_ ( .A1(\myexu/myalu/_0601_ ), .A2(\myexu/myalu/_1363_ ), .ZN(\myexu/myalu/_0606_ ) );
NOR3_X1 \myexu/myalu/_1588_ ( .A1(\myexu/myalu/_1364_ ), .A2(\myexu/myalu/_1365_ ), .A3(\myexu/myalu/_1366_ ), .ZN(\myexu/myalu/_0607_ ) );
NOR2_X1 \myexu/myalu/_1589_ ( .A1(\myexu/myalu/_1367_ ), .A2(\myexu/myalu/_1368_ ), .ZN(\myexu/myalu/_0608_ ) );
INV_X1 \myexu/myalu/_1590_ ( .A(\myexu/myalu/_1369_ ), .ZN(\myexu/myalu/_0609_ ) );
AND3_X1 \myexu/myalu/_1591_ ( .A1(\myexu/myalu/_0608_ ), .A2(\myexu/myalu/_0609_ ), .A3(\myexu/myalu/_0539_ ), .ZN(\myexu/myalu/_0610_ ) );
NOR2_X1 \myexu/myalu/_1592_ ( .A1(\myexu/myalu/_1372_ ), .A2(\myexu/myalu/_1373_ ), .ZN(\myexu/myalu/_0611_ ) );
NOR2_X1 \myexu/myalu/_1593_ ( .A1(\myexu/myalu/_1374_ ), .A2(\myexu/myalu/_1375_ ), .ZN(\myexu/myalu/_0612_ ) );
AND3_X1 \myexu/myalu/_1594_ ( .A1(\myexu/myalu/_0610_ ), .A2(\myexu/myalu/_0611_ ), .A3(\myexu/myalu/_0612_ ), .ZN(\myexu/myalu/_0613_ ) );
NOR2_X1 \myexu/myalu/_1595_ ( .A1(\myexu/myalu/_1378_ ), .A2(\myexu/myalu/_1379_ ), .ZN(\myexu/myalu/_0614_ ) );
AND3_X1 \myexu/myalu/_1596_ ( .A1(\myexu/myalu/_0614_ ), .A2(\myexu/myalu/_0561_ ), .A3(\myexu/myalu/_0563_ ), .ZN(\myexu/myalu/_0615_ ) );
NOR2_X1 \myexu/myalu/_1597_ ( .A1(\myexu/myalu/_1380_ ), .A2(\myexu/myalu/_1381_ ), .ZN(\myexu/myalu/_0616_ ) );
AND3_X1 \myexu/myalu/_1598_ ( .A1(\myexu/myalu/_0616_ ), .A2(\myexu/myalu/_0557_ ), .A3(\myexu/myalu/_0573_ ), .ZN(\myexu/myalu/_0617_ ) );
AND2_X1 \myexu/myalu/_1599_ ( .A1(\myexu/myalu/_0615_ ), .A2(\myexu/myalu/_0617_ ), .ZN(\myexu/myalu/_0618_ ) );
NAND2_X1 \myexu/myalu/_1600_ ( .A1(\myexu/myalu/_0613_ ), .A2(\myexu/myalu/_0618_ ), .ZN(\myexu/myalu/_0619_ ) );
NAND3_X1 \myexu/myalu/_1601_ ( .A1(\myexu/myalu/_0606_ ), .A2(\myexu/myalu/_0607_ ), .A3(\myexu/myalu/_0619_ ), .ZN(\myexu/myalu/_0620_ ) );
NAND2_X1 \myexu/myalu/_1602_ ( .A1(\myexu/myalu/_0605_ ), .A2(\myexu/myalu/_0620_ ), .ZN(\myexu/myalu/_0621_ ) );
AND2_X1 \myexu/myalu/_1603_ ( .A1(\myexu/myalu/_1372_ ), .A2(\myexu/myalu/_1373_ ), .ZN(\myexu/myalu/_0622_ ) );
AND3_X1 \myexu/myalu/_1604_ ( .A1(\myexu/myalu/_0622_ ), .A2(\myexu/myalu/_1374_ ), .A3(\myexu/myalu/_1375_ ), .ZN(\myexu/myalu/_0623_ ) );
AND2_X1 \myexu/myalu/_1605_ ( .A1(\myexu/myalu/_1383_ ), .A2(\myexu/myalu/_1384_ ), .ZN(\myexu/myalu/_0624_ ) );
AND3_X1 \myexu/myalu/_1606_ ( .A1(\myexu/myalu/_0624_ ), .A2(\myexu/myalu/_1380_ ), .A3(\myexu/myalu/_1381_ ), .ZN(\myexu/myalu/_0625_ ) );
AND4_X1 \myexu/myalu/_1607_ ( .A1(\myexu/myalu/_1376_ ), .A2(\myexu/myalu/_1377_ ), .A3(\myexu/myalu/_1378_ ), .A4(\myexu/myalu/_1379_ ), .ZN(\myexu/myalu/_0626_ ) );
AND3_X1 \myexu/myalu/_1608_ ( .A1(\myexu/myalu/_0623_ ), .A2(\myexu/myalu/_0625_ ), .A3(\myexu/myalu/_0626_ ), .ZN(\myexu/myalu/_0627_ ) );
AND4_X1 \myexu/myalu/_1609_ ( .A1(\myexu/myalu/_1367_ ), .A2(\myexu/myalu/_1368_ ), .A3(\myexu/myalu/_1369_ ), .A4(\myexu/myalu/_1370_ ), .ZN(\myexu/myalu/_0628_ ) );
AND4_X1 \myexu/myalu/_1610_ ( .A1(\myexu/myalu/_1363_ ), .A2(\myexu/myalu/_1364_ ), .A3(\myexu/myalu/_1365_ ), .A4(\myexu/myalu/_1366_ ), .ZN(\myexu/myalu/_0629_ ) );
NAND3_X1 \myexu/myalu/_1611_ ( .A1(\myexu/myalu/_0627_ ), .A2(\myexu/myalu/_0628_ ), .A3(\myexu/myalu/_0629_ ), .ZN(\myexu/myalu/_0630_ ) );
AOI21_X1 \myexu/myalu/_1612_ ( .A(\myexu/myalu/_0630_ ), .B1(\myexu/myalu/_0598_ ), .B2(\myexu/myalu/_0599_ ), .ZN(\myexu/myalu/_0631_ ) );
AOI21_X1 \myexu/myalu/_1613_ ( .A(\myexu/myalu/_0631_ ), .B1(\myexu/myalu/_0606_ ), .B2(\myexu/myalu/_0607_ ), .ZN(\myexu/myalu/_0632_ ) );
NOR2_X4 \myexu/myalu/_1614_ ( .A1(\myexu/myalu/_0621_ ), .A2(\myexu/myalu/_0632_ ), .ZN(\myexu/myalu/_0633_ ) );
BUF_X4 \myexu/myalu/_1615_ ( .A(\myexu/myalu/_0633_ ), .Z(\myexu/myalu/_0634_ ) );
AND2_X2 \myexu/myalu/_1616_ ( .A1(\myexu/myalu/_0001_ ), .A2(\myexu/myalu/_0000_ ), .ZN(\myexu/myalu/_0635_ ) );
AND2_X2 \myexu/myalu/_1617_ ( .A1(\myexu/myalu/_0635_ ), .A2(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0636_ ) );
AND4_X1 \myexu/myalu/_1618_ ( .A1(\myexu/myalu/_1387_ ), .A2(\myexu/myalu/_0634_ ), .A3(\myexu/myalu/_0589_ ), .A4(\myexu/myalu/_0636_ ), .ZN(\myexu/myalu/_0637_ ) );
NOR2_X1 \myexu/myalu/_1619_ ( .A1(\myexu/myalu/_0515_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0638_ ) );
AND2_X1 \myexu/myalu/_1620_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1330_ ), .ZN(\myexu/myalu/_0639_ ) );
INV_X1 \myexu/myalu/_1621_ ( .A(fanout_net_11 ), .ZN(\myexu/myalu/_0640_ ) );
BUF_X2 \myexu/myalu/_1622_ ( .A(\myexu/myalu/_0640_ ), .Z(\myexu/myalu/_0641_ ) );
OR3_X1 \myexu/myalu/_1623_ ( .A1(\myexu/myalu/_0638_ ), .A2(\myexu/myalu/_0639_ ), .A3(\myexu/myalu/_0641_ ), .ZN(\myexu/myalu/_0642_ ) );
NOR2_X1 \myexu/myalu/_1624_ ( .A1(\myexu/myalu/_0510_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0643_ ) );
AND2_X1 \myexu/myalu/_1625_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1359_ ), .ZN(\myexu/myalu/_0644_ ) );
OR3_X1 \myexu/myalu/_1626_ ( .A1(\myexu/myalu/_0643_ ), .A2(\myexu/myalu/_0644_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0645_ ) );
BUF_X4 \myexu/myalu/_1627_ ( .A(\myexu/myalu/_0585_ ), .Z(\myexu/myalu/_0646_ ) );
NAND3_X1 \myexu/myalu/_1628_ ( .A1(\myexu/myalu/_0642_ ), .A2(\myexu/myalu/_0645_ ), .A3(\myexu/myalu/_0646_ ), .ZN(\myexu/myalu/_0647_ ) );
NOR2_X1 \myexu/myalu/_1629_ ( .A1(\myexu/myalu/_0526_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0648_ ) );
AND2_X1 \myexu/myalu/_1630_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1334_ ), .ZN(\myexu/myalu/_0649_ ) );
OR3_X1 \myexu/myalu/_1631_ ( .A1(\myexu/myalu/_0648_ ), .A2(\myexu/myalu/_0649_ ), .A3(\myexu/myalu/_0640_ ), .ZN(\myexu/myalu/_0650_ ) );
NOR2_X1 \myexu/myalu/_1632_ ( .A1(\myexu/myalu/_0521_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0651_ ) );
AND2_X1 \myexu/myalu/_1633_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1332_ ), .ZN(\myexu/myalu/_0652_ ) );
OR3_X1 \myexu/myalu/_1634_ ( .A1(\myexu/myalu/_0651_ ), .A2(\myexu/myalu/_0652_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0653_ ) );
NAND3_X1 \myexu/myalu/_1635_ ( .A1(\myexu/myalu/_0650_ ), .A2(\myexu/myalu/_0653_ ), .A3(fanout_net_13 ), .ZN(\myexu/myalu/_0654_ ) );
AOI21_X1 \myexu/myalu/_1636_ ( .A(\myexu/myalu/_0505_ ), .B1(\myexu/myalu/_0647_ ), .B2(\myexu/myalu/_0654_ ), .ZN(\myexu/myalu/_0655_ ) );
NAND2_X1 \myexu/myalu/_1637_ ( .A1(\myexu/myalu/_0584_ ), .A2(\myexu/myalu/_1328_ ), .ZN(\myexu/myalu/_0656_ ) );
INV_X1 \myexu/myalu/_1638_ ( .A(fanout_net_9 ), .ZN(\myexu/myalu/_0657_ ) );
BUF_X2 \myexu/myalu/_1639_ ( .A(\myexu/myalu/_0657_ ), .Z(\myexu/myalu/_0658_ ) );
NOR2_X1 \myexu/myalu/_1640_ ( .A1(\myexu/myalu/_0658_ ), .A2(fanout_net_11 ), .ZN(\myexu/myalu/_0659_ ) );
INV_X1 \myexu/myalu/_1641_ ( .A(\myexu/myalu/_0659_ ), .ZN(\myexu/myalu/_0660_ ) );
NOR2_X1 \myexu/myalu/_1642_ ( .A1(\myexu/myalu/_0502_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0661_ ) );
AND2_X1 \myexu/myalu/_1643_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1353_ ), .ZN(\myexu/myalu/_0662_ ) );
NOR2_X1 \myexu/myalu/_1644_ ( .A1(\myexu/myalu/_0661_ ), .A2(\myexu/myalu/_0662_ ), .ZN(\myexu/myalu/_0663_ ) );
BUF_X2 \myexu/myalu/_1645_ ( .A(\myexu/myalu/_0640_ ), .Z(\myexu/myalu/_0664_ ) );
OAI221_X1 \myexu/myalu/_1646_ ( .A(\myexu/myalu/_0656_ ), .B1(\myexu/myalu/_0660_ ), .B2(\myexu/myalu/_0499_ ), .C1(\myexu/myalu/_0663_ ), .C2(\myexu/myalu/_0664_ ), .ZN(\myexu/myalu/_0665_ ) );
NOR2_X1 \myexu/myalu/_1647_ ( .A1(\myexu/myalu/_0476_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0666_ ) );
AND2_X1 \myexu/myalu/_1648_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1357_ ), .ZN(\myexu/myalu/_0667_ ) );
OR3_X1 \myexu/myalu/_1649_ ( .A1(\myexu/myalu/_0666_ ), .A2(\myexu/myalu/_0667_ ), .A3(\myexu/myalu/_0640_ ), .ZN(\myexu/myalu/_0668_ ) );
NOR2_X1 \myexu/myalu/_1650_ ( .A1(\myexu/myalu/_0483_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0669_ ) );
AND2_X1 \myexu/myalu/_1651_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1355_ ), .ZN(\myexu/myalu/_0670_ ) );
OR3_X1 \myexu/myalu/_1652_ ( .A1(\myexu/myalu/_0669_ ), .A2(\myexu/myalu/_0670_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0671_ ) );
AND2_X1 \myexu/myalu/_1653_ ( .A1(\myexu/myalu/_0668_ ), .A2(\myexu/myalu/_0671_ ), .ZN(\myexu/myalu/_0672_ ) );
MUX2_X1 \myexu/myalu/_1654_ ( .A(\myexu/myalu/_0665_ ), .B(\myexu/myalu/_0672_ ), .S(fanout_net_13 ), .Z(\myexu/myalu/_0673_ ) );
AOI211_X4 \myexu/myalu/_1655_ ( .A(fanout_net_17 ), .B(\myexu/myalu/_0655_ ), .C1(\myexu/myalu/_0673_ ), .C2(\myexu/myalu/_0506_ ), .ZN(\myexu/myalu/_0674_ ) );
INV_X1 \myexu/myalu/_1656_ ( .A(\myexu/myalu/_0001_ ), .ZN(\myexu/myalu/_0675_ ) );
NOR2_X2 \myexu/myalu/_1657_ ( .A1(\myexu/myalu/_0675_ ), .A2(\myexu/myalu/_0000_ ), .ZN(\myexu/myalu/_0676_ ) );
AND2_X1 \myexu/myalu/_1658_ ( .A1(\myexu/myalu/_0676_ ), .A2(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0677_ ) );
NOR2_X1 \myexu/myalu/_1659_ ( .A1(\myexu/myalu/_0677_ ), .A2(\myexu/myalu/_0636_ ), .ZN(\myexu/myalu/_0678_ ) );
NOR2_X1 \myexu/myalu/_1660_ ( .A1(\myexu/myalu/_0566_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0679_ ) );
AND2_X1 \myexu/myalu/_1661_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1347_ ), .ZN(\myexu/myalu/_0680_ ) );
OR3_X1 \myexu/myalu/_1662_ ( .A1(\myexu/myalu/_0679_ ), .A2(\myexu/myalu/_0680_ ), .A3(\myexu/myalu/_0640_ ), .ZN(\myexu/myalu/_0681_ ) );
INV_X1 \myexu/myalu/_1663_ ( .A(\myexu/myalu/_1344_ ), .ZN(\myexu/myalu/_0682_ ) );
NOR2_X1 \myexu/myalu/_1664_ ( .A1(\myexu/myalu/_0682_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0683_ ) );
AND2_X1 \myexu/myalu/_1665_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1345_ ), .ZN(\myexu/myalu/_0684_ ) );
OR3_X1 \myexu/myalu/_1666_ ( .A1(\myexu/myalu/_0683_ ), .A2(\myexu/myalu/_0684_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0685_ ) );
AND2_X1 \myexu/myalu/_1667_ ( .A1(\myexu/myalu/_0681_ ), .A2(\myexu/myalu/_0685_ ), .ZN(\myexu/myalu/_0686_ ) );
MUX2_X1 \myexu/myalu/_1668_ ( .A(\myexu/myalu/_1351_ ), .B(\myexu/myalu/_1352_ ), .S(fanout_net_9 ), .Z(\myexu/myalu/_0687_ ) );
OR2_X1 \myexu/myalu/_1669_ ( .A1(\myexu/myalu/_0687_ ), .A2(\myexu/myalu/_0640_ ), .ZN(\myexu/myalu/_0688_ ) );
NOR2_X1 \myexu/myalu/_1670_ ( .A1(\myexu/myalu/_0575_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0689_ ) );
AND2_X1 \myexu/myalu/_1671_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1349_ ), .ZN(\myexu/myalu/_0690_ ) );
OR3_X1 \myexu/myalu/_1672_ ( .A1(\myexu/myalu/_0689_ ), .A2(\myexu/myalu/_0690_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0691_ ) );
AND2_X1 \myexu/myalu/_1673_ ( .A1(\myexu/myalu/_0688_ ), .A2(\myexu/myalu/_0691_ ), .ZN(\myexu/myalu/_0692_ ) );
MUX2_X1 \myexu/myalu/_1674_ ( .A(\myexu/myalu/_0686_ ), .B(\myexu/myalu/_0692_ ), .S(fanout_net_13 ), .Z(\myexu/myalu/_0693_ ) );
OR2_X1 \myexu/myalu/_1675_ ( .A1(\myexu/myalu/_0693_ ), .A2(\myexu/myalu/_0506_ ), .ZN(\myexu/myalu/_0694_ ) );
BUF_X2 \myexu/myalu/_1676_ ( .A(\myexu/myalu/_0664_ ), .Z(\myexu/myalu/_0695_ ) );
NOR2_X1 \myexu/myalu/_1677_ ( .A1(\myexu/myalu/_0534_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0696_ ) );
AND2_X1 \myexu/myalu/_1678_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1336_ ), .ZN(\myexu/myalu/_0697_ ) );
OAI21_X1 \myexu/myalu/_1679_ ( .A(\myexu/myalu/_0695_ ), .B1(\myexu/myalu/_0696_ ), .B2(\myexu/myalu/_0697_ ), .ZN(\myexu/myalu/_0698_ ) );
NOR2_X1 \myexu/myalu/_1680_ ( .A1(\myexu/myalu/_0542_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0699_ ) );
AND2_X1 \myexu/myalu/_1681_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1338_ ), .ZN(\myexu/myalu/_0700_ ) );
OAI21_X1 \myexu/myalu/_1682_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0699_ ), .B2(\myexu/myalu/_0700_ ), .ZN(\myexu/myalu/_0701_ ) );
NAND2_X1 \myexu/myalu/_1683_ ( .A1(\myexu/myalu/_0698_ ), .A2(\myexu/myalu/_0701_ ), .ZN(\myexu/myalu/_0702_ ) );
BUF_X4 \myexu/myalu/_1684_ ( .A(\myexu/myalu/_0646_ ), .Z(\myexu/myalu/_0703_ ) );
NAND2_X1 \myexu/myalu/_1685_ ( .A1(\myexu/myalu/_0702_ ), .A2(\myexu/myalu/_0703_ ), .ZN(\myexu/myalu/_0704_ ) );
NOR2_X1 \myexu/myalu/_1686_ ( .A1(\myexu/myalu/_0549_ ), .A2(fanout_net_9 ), .ZN(\myexu/myalu/_0705_ ) );
AND2_X1 \myexu/myalu/_1687_ ( .A1(fanout_net_9 ), .A2(\myexu/myalu/_1341_ ), .ZN(\myexu/myalu/_0706_ ) );
OAI21_X1 \myexu/myalu/_1688_ ( .A(\myexu/myalu/_0641_ ), .B1(\myexu/myalu/_0705_ ), .B2(\myexu/myalu/_0706_ ), .ZN(\myexu/myalu/_0707_ ) );
NOR2_X1 \myexu/myalu/_1689_ ( .A1(\myexu/myalu/_0545_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0708_ ) );
AND2_X1 \myexu/myalu/_1690_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1343_ ), .ZN(\myexu/myalu/_0709_ ) );
OAI21_X1 \myexu/myalu/_1691_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0708_ ), .B2(\myexu/myalu/_0709_ ), .ZN(\myexu/myalu/_0710_ ) );
NAND2_X1 \myexu/myalu/_1692_ ( .A1(\myexu/myalu/_0707_ ), .A2(\myexu/myalu/_0710_ ), .ZN(\myexu/myalu/_0711_ ) );
NAND2_X1 \myexu/myalu/_1693_ ( .A1(\myexu/myalu/_0711_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0712_ ) );
NAND2_X1 \myexu/myalu/_1694_ ( .A1(\myexu/myalu/_0704_ ), .A2(\myexu/myalu/_0712_ ), .ZN(\myexu/myalu/_0713_ ) );
OAI21_X1 \myexu/myalu/_1695_ ( .A(\myexu/myalu/_0694_ ), .B1(fanout_net_15 ), .B2(\myexu/myalu/_0713_ ), .ZN(\myexu/myalu/_0714_ ) );
AOI211_X4 \myexu/myalu/_1696_ ( .A(\myexu/myalu/_0674_ ), .B(\myexu/myalu/_0678_ ), .C1(\myexu/myalu/_0714_ ), .C2(fanout_net_17 ), .ZN(\myexu/myalu/_0715_ ) );
AND2_X1 \myexu/myalu/_1697_ ( .A1(\myexu/myalu/_0675_ ), .A2(\myexu/myalu/_0000_ ), .ZN(\myexu/myalu/_0716_ ) );
AND2_X1 \myexu/myalu/_1698_ ( .A1(\myexu/myalu/_0716_ ), .A2(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0717_ ) );
AND2_X1 \myexu/myalu/_1699_ ( .A1(\myexu/myalu/_0717_ ), .A2(\myexu/myalu/_0588_ ), .ZN(\myexu/myalu/_0718_ ) );
AND3_X1 \myexu/myalu/_1700_ ( .A1(\myexu/myalu/_0718_ ), .A2(\myexu/myalu/_1328_ ), .A3(\myexu/myalu/_0587_ ), .ZN(\myexu/myalu/_0719_ ) );
XNOR2_X1 \myexu/myalu/_1701_ ( .A(fanout_net_10 ), .B(\myexu/myalu/_1328_ ), .ZN(\myexu/myalu/_0720_ ) );
AND2_X2 \myexu/myalu/_1702_ ( .A1(\myexu/myalu/_0635_ ), .A2(\myexu/myalu/_0572_ ), .ZN(\myexu/myalu/_0721_ ) );
INV_X1 \myexu/myalu/_1703_ ( .A(\myexu/myalu/_0721_ ), .ZN(\myexu/myalu/_0722_ ) );
AND2_X1 \myexu/myalu/_1704_ ( .A1(\myexu/myalu/_0559_ ), .A2(\myexu/myalu/_0572_ ), .ZN(\myexu/myalu/_0723_ ) );
INV_X1 \myexu/myalu/_1705_ ( .A(\myexu/myalu/_0723_ ), .ZN(\myexu/myalu/_0724_ ) );
AOI21_X1 \myexu/myalu/_1706_ ( .A(\myexu/myalu/_0720_ ), .B1(\myexu/myalu/_0722_ ), .B2(\myexu/myalu/_0724_ ), .ZN(\myexu/myalu/_0725_ ) );
AND2_X2 \myexu/myalu/_1707_ ( .A1(\myexu/myalu/_0676_ ), .A2(\myexu/myalu/_0572_ ), .ZN(\myexu/myalu/_0726_ ) );
OAI21_X1 \myexu/myalu/_1708_ ( .A(\myexu/myalu/_0726_ ), .B1(fanout_net_10 ), .B2(\myexu/myalu/_1328_ ), .ZN(\myexu/myalu/_0727_ ) );
BUF_X4 \myexu/myalu/_1709_ ( .A(\myexu/myalu/_0716_ ), .Z(\myexu/myalu/_0728_ ) );
BUF_X4 \myexu/myalu/_1710_ ( .A(\myexu/myalu/_0572_ ), .Z(\myexu/myalu/_0729_ ) );
AND2_X1 \myexu/myalu/_1711_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1328_ ), .ZN(\myexu/myalu/_0730_ ) );
NAND3_X1 \myexu/myalu/_1712_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0729_ ), .A3(\myexu/myalu/_0730_ ), .ZN(\myexu/myalu/_0731_ ) );
NAND2_X1 \myexu/myalu/_1713_ ( .A1(\myexu/myalu/_0727_ ), .A2(\myexu/myalu/_0731_ ), .ZN(\myexu/myalu/_0732_ ) );
OR3_X1 \myexu/myalu/_1714_ ( .A1(\myexu/myalu/_0719_ ), .A2(\myexu/myalu/_0725_ ), .A3(\myexu/myalu/_0732_ ), .ZN(\myexu/myalu/_0733_ ) );
OR4_X1 \myexu/myalu/_1715_ ( .A1(\myexu/myalu/_0581_ ), .A2(\myexu/myalu/_0637_ ), .A3(\myexu/myalu/_0715_ ), .A4(\myexu/myalu/_0733_ ), .ZN(\myexu/myalu/_1296_ ) );
INV_X1 \myexu/myalu/_1716_ ( .A(\myexu/myalu/_0677_ ), .ZN(\myexu/myalu/_0734_ ) );
AND2_X1 \myexu/myalu/_1717_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_1338_ ), .ZN(\myexu/myalu/_0735_ ) );
AND2_X1 \myexu/myalu/_1718_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1340_ ), .ZN(\myexu/myalu/_0736_ ) );
OAI21_X1 \myexu/myalu/_1719_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0735_ ), .B2(\myexu/myalu/_0736_ ), .ZN(\myexu/myalu/_0737_ ) );
NOR2_X1 \myexu/myalu/_1720_ ( .A1(\myexu/myalu/_0536_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0738_ ) );
AND2_X1 \myexu/myalu/_1721_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1337_ ), .ZN(\myexu/myalu/_0739_ ) );
OAI21_X1 \myexu/myalu/_1722_ ( .A(\myexu/myalu/_0641_ ), .B1(\myexu/myalu/_0738_ ), .B2(\myexu/myalu/_0739_ ), .ZN(\myexu/myalu/_0740_ ) );
NAND2_X1 \myexu/myalu/_1723_ ( .A1(\myexu/myalu/_0737_ ), .A2(\myexu/myalu/_0740_ ), .ZN(\myexu/myalu/_0741_ ) );
NAND2_X1 \myexu/myalu/_1724_ ( .A1(\myexu/myalu/_0741_ ), .A2(\myexu/myalu/_0646_ ), .ZN(\myexu/myalu/_0742_ ) );
AND2_X1 \myexu/myalu/_1725_ ( .A1(\myexu/myalu/_0657_ ), .A2(\myexu/myalu/_1343_ ), .ZN(\myexu/myalu/_0743_ ) );
AND2_X1 \myexu/myalu/_1726_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1344_ ), .ZN(\myexu/myalu/_0744_ ) );
OAI21_X1 \myexu/myalu/_1727_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0743_ ), .B2(\myexu/myalu/_0744_ ), .ZN(\myexu/myalu/_0745_ ) );
NOR2_X1 \myexu/myalu/_1728_ ( .A1(\myexu/myalu/_0551_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0746_ ) );
AND2_X1 \myexu/myalu/_1729_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1342_ ), .ZN(\myexu/myalu/_0747_ ) );
OAI21_X1 \myexu/myalu/_1730_ ( .A(\myexu/myalu/_0641_ ), .B1(\myexu/myalu/_0746_ ), .B2(\myexu/myalu/_0747_ ), .ZN(\myexu/myalu/_0748_ ) );
NAND2_X1 \myexu/myalu/_1731_ ( .A1(\myexu/myalu/_0745_ ), .A2(\myexu/myalu/_0748_ ), .ZN(\myexu/myalu/_0749_ ) );
NAND2_X1 \myexu/myalu/_1732_ ( .A1(\myexu/myalu/_0749_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0750_ ) );
NAND2_X1 \myexu/myalu/_1733_ ( .A1(\myexu/myalu/_0742_ ), .A2(\myexu/myalu/_0750_ ), .ZN(\myexu/myalu/_0751_ ) );
NAND3_X1 \myexu/myalu/_1734_ ( .A1(\myexu/myalu/_0658_ ), .A2(fanout_net_11 ), .A3(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_0752_ ) );
INV_X1 \myexu/myalu/_1735_ ( .A(\myexu/myalu/_1351_ ), .ZN(\myexu/myalu/_0753_ ) );
MUX2_X1 \myexu/myalu/_1736_ ( .A(\myexu/myalu/_0577_ ), .B(\myexu/myalu/_0753_ ), .S(fanout_net_10 ), .Z(\myexu/myalu/_0754_ ) );
OAI21_X1 \myexu/myalu/_1737_ ( .A(\myexu/myalu/_0752_ ), .B1(\myexu/myalu/_0754_ ), .B2(fanout_net_11 ), .ZN(\myexu/myalu/_0755_ ) );
AND2_X1 \myexu/myalu/_1738_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_1345_ ), .ZN(\myexu/myalu/_0756_ ) );
AND2_X1 \myexu/myalu/_1739_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1346_ ), .ZN(\myexu/myalu/_0757_ ) );
OAI21_X1 \myexu/myalu/_1740_ ( .A(\myexu/myalu/_0641_ ), .B1(\myexu/myalu/_0756_ ), .B2(\myexu/myalu/_0757_ ), .ZN(\myexu/myalu/_0758_ ) );
NOR2_X1 \myexu/myalu/_1741_ ( .A1(\myexu/myalu/_0568_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0759_ ) );
AND2_X1 \myexu/myalu/_1742_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1348_ ), .ZN(\myexu/myalu/_0760_ ) );
OAI21_X1 \myexu/myalu/_1743_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0759_ ), .B2(\myexu/myalu/_0760_ ), .ZN(\myexu/myalu/_0761_ ) );
NAND2_X1 \myexu/myalu/_1744_ ( .A1(\myexu/myalu/_0758_ ), .A2(\myexu/myalu/_0761_ ), .ZN(\myexu/myalu/_0762_ ) );
MUX2_X1 \myexu/myalu/_1745_ ( .A(\myexu/myalu/_0755_ ), .B(\myexu/myalu/_0762_ ), .S(\myexu/myalu/_0646_ ), .Z(\myexu/myalu/_0763_ ) );
MUX2_X1 \myexu/myalu/_1746_ ( .A(\myexu/myalu/_0751_ ), .B(\myexu/myalu/_0763_ ), .S(fanout_net_15 ), .Z(\myexu/myalu/_0764_ ) );
NAND2_X1 \myexu/myalu/_1747_ ( .A1(\myexu/myalu/_0764_ ), .A2(fanout_net_17 ), .ZN(\myexu/myalu/_0765_ ) );
AND2_X1 \myexu/myalu/_1748_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_1330_ ), .ZN(\myexu/myalu/_0766_ ) );
AND2_X1 \myexu/myalu/_1749_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1331_ ), .ZN(\myexu/myalu/_0767_ ) );
OAI21_X1 \myexu/myalu/_1750_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0766_ ), .B2(\myexu/myalu/_0767_ ), .ZN(\myexu/myalu/_0768_ ) );
NOR2_X1 \myexu/myalu/_1751_ ( .A1(\myexu/myalu/_0512_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0769_ ) );
AND2_X1 \myexu/myalu/_1752_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1329_ ), .ZN(\myexu/myalu/_0770_ ) );
OAI21_X1 \myexu/myalu/_1753_ ( .A(\myexu/myalu/_0664_ ), .B1(\myexu/myalu/_0769_ ), .B2(\myexu/myalu/_0770_ ), .ZN(\myexu/myalu/_0771_ ) );
NAND2_X1 \myexu/myalu/_1754_ ( .A1(\myexu/myalu/_0768_ ), .A2(\myexu/myalu/_0771_ ), .ZN(\myexu/myalu/_0772_ ) );
BUF_X2 \myexu/myalu/_1755_ ( .A(\myexu/myalu/_0646_ ), .Z(\myexu/myalu/_0773_ ) );
NAND2_X1 \myexu/myalu/_1756_ ( .A1(\myexu/myalu/_0772_ ), .A2(\myexu/myalu/_0773_ ), .ZN(\myexu/myalu/_0774_ ) );
AND2_X1 \myexu/myalu/_1757_ ( .A1(\myexu/myalu/_0657_ ), .A2(\myexu/myalu/_1334_ ), .ZN(\myexu/myalu/_0775_ ) );
AND2_X1 \myexu/myalu/_1758_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1335_ ), .ZN(\myexu/myalu/_0776_ ) );
OR3_X1 \myexu/myalu/_1759_ ( .A1(\myexu/myalu/_0775_ ), .A2(\myexu/myalu/_0640_ ), .A3(\myexu/myalu/_0776_ ), .ZN(\myexu/myalu/_0777_ ) );
NOR2_X1 \myexu/myalu/_1760_ ( .A1(\myexu/myalu/_0523_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0778_ ) );
AND2_X1 \myexu/myalu/_1761_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1333_ ), .ZN(\myexu/myalu/_0779_ ) );
OR3_X1 \myexu/myalu/_1762_ ( .A1(\myexu/myalu/_0778_ ), .A2(\myexu/myalu/_0779_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0780_ ) );
NAND3_X1 \myexu/myalu/_1763_ ( .A1(\myexu/myalu/_0777_ ), .A2(fanout_net_13 ), .A3(\myexu/myalu/_0780_ ), .ZN(\myexu/myalu/_0781_ ) );
AND3_X1 \myexu/myalu/_1764_ ( .A1(\myexu/myalu/_0774_ ), .A2(\myexu/myalu/_0781_ ), .A3(fanout_net_15 ), .ZN(\myexu/myalu/_0782_ ) );
AND2_X1 \myexu/myalu/_1765_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_1353_ ), .ZN(\myexu/myalu/_0783_ ) );
AND2_X1 \myexu/myalu/_1766_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1354_ ), .ZN(\myexu/myalu/_0784_ ) );
OAI21_X1 \myexu/myalu/_1767_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0783_ ), .B2(\myexu/myalu/_0784_ ), .ZN(\myexu/myalu/_0785_ ) );
MUX2_X1 \myexu/myalu/_1768_ ( .A(\myexu/myalu/_0499_ ), .B(\myexu/myalu/_0502_ ), .S(fanout_net_10 ), .Z(\myexu/myalu/_0786_ ) );
OAI211_X2 \myexu/myalu/_1769_ ( .A(\myexu/myalu/_0785_ ), .B(\myexu/myalu/_0773_ ), .C1(fanout_net_11 ), .C2(\myexu/myalu/_0786_ ), .ZN(\myexu/myalu/_0787_ ) );
BUF_X4 \myexu/myalu/_1770_ ( .A(\myexu/myalu/_0641_ ), .Z(\myexu/myalu/_0788_ ) );
AND2_X1 \myexu/myalu/_1771_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_1355_ ), .ZN(\myexu/myalu/_0789_ ) );
AND2_X1 \myexu/myalu/_1772_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1356_ ), .ZN(\myexu/myalu/_0790_ ) );
OAI21_X1 \myexu/myalu/_1773_ ( .A(\myexu/myalu/_0788_ ), .B1(\myexu/myalu/_0789_ ), .B2(\myexu/myalu/_0790_ ), .ZN(\myexu/myalu/_0791_ ) );
NOR2_X1 \myexu/myalu/_1774_ ( .A1(\myexu/myalu/_0481_ ), .A2(fanout_net_10 ), .ZN(\myexu/myalu/_0792_ ) );
AND2_X1 \myexu/myalu/_1775_ ( .A1(fanout_net_10 ), .A2(\myexu/myalu/_1358_ ), .ZN(\myexu/myalu/_0793_ ) );
OAI21_X1 \myexu/myalu/_1776_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0792_ ), .B2(\myexu/myalu/_0793_ ), .ZN(\myexu/myalu/_0794_ ) );
NAND3_X1 \myexu/myalu/_1777_ ( .A1(\myexu/myalu/_0791_ ), .A2(fanout_net_13 ), .A3(\myexu/myalu/_0794_ ), .ZN(\myexu/myalu/_0795_ ) );
AOI21_X1 \myexu/myalu/_1778_ ( .A(fanout_net_15 ), .B1(\myexu/myalu/_0787_ ), .B2(\myexu/myalu/_0795_ ), .ZN(\myexu/myalu/_0796_ ) );
OR3_X1 \myexu/myalu/_1779_ ( .A1(\myexu/myalu/_0782_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0796_ ), .ZN(\myexu/myalu/_0797_ ) );
AOI21_X1 \myexu/myalu/_1780_ ( .A(\myexu/myalu/_0734_ ), .B1(\myexu/myalu/_0765_ ), .B2(\myexu/myalu/_0797_ ), .ZN(\myexu/myalu/_0798_ ) );
MUX2_X1 \myexu/myalu/_1781_ ( .A(\myexu/myalu/_0499_ ), .B(\myexu/myalu/_0497_ ), .S(fanout_net_10 ), .Z(\myexu/myalu/_0799_ ) );
OR3_X1 \myexu/myalu/_1782_ ( .A1(\myexu/myalu/_0799_ ), .A2(fanout_net_13 ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0800_ ) );
INV_X1 \myexu/myalu/_1783_ ( .A(\myexu/myalu/_0717_ ), .ZN(\myexu/myalu/_0801_ ) );
NOR4_X1 \myexu/myalu/_1784_ ( .A1(\myexu/myalu/_0800_ ), .A2(\myexu/myalu/_0801_ ), .A3(fanout_net_17 ), .A4(fanout_net_15 ), .ZN(\myexu/myalu/_0802_ ) );
XNOR2_X1 \myexu/myalu/_1785_ ( .A(\myexu/myalu/_0586_ ), .B(\myexu/myalu/_0505_ ), .ZN(\myexu/myalu/_0803_ ) );
NOR2_X1 \myexu/myalu/_1786_ ( .A1(\myexu/myalu/_0584_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0804_ ) );
INV_X1 \myexu/myalu/_1787_ ( .A(\myexu/myalu/_0804_ ), .ZN(\myexu/myalu/_0805_ ) );
NAND3_X1 \myexu/myalu/_1788_ ( .A1(\myexu/myalu/_0633_ ), .A2(\myexu/myalu/_0803_ ), .A3(\myexu/myalu/_0805_ ), .ZN(\myexu/myalu/_0806_ ) );
NOR3_X1 \myexu/myalu/_1789_ ( .A1(\myexu/myalu/_0585_ ), .A2(fanout_net_10 ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0807_ ) );
NOR2_X2 \myexu/myalu/_1790_ ( .A1(\myexu/myalu/_0806_ ), .A2(\myexu/myalu/_0807_ ), .ZN(\myexu/myalu/_0808_ ) );
XNOR2_X1 \myexu/myalu/_1791_ ( .A(fanout_net_10 ), .B(fanout_net_11 ), .ZN(\myexu/myalu/_0809_ ) );
XNOR2_X1 \myexu/myalu/_1792_ ( .A(\myexu/myalu/_0589_ ), .B(\myexu/myalu/_1387_ ), .ZN(\myexu/myalu/_0810_ ) );
XNOR2_X1 \myexu/myalu/_1793_ ( .A(\myexu/myalu/_0587_ ), .B(\myexu/myalu/_0588_ ), .ZN(\myexu/myalu/_0811_ ) );
AND2_X2 \myexu/myalu/_1794_ ( .A1(\myexu/myalu/_0810_ ), .A2(\myexu/myalu/_0811_ ), .ZN(\myexu/myalu/_0812_ ) );
NAND3_X1 \myexu/myalu/_1795_ ( .A1(\myexu/myalu/_0808_ ), .A2(\myexu/myalu/_0809_ ), .A3(\myexu/myalu/_0812_ ), .ZN(\myexu/myalu/_0813_ ) );
NAND3_X1 \myexu/myalu/_1796_ ( .A1(\myexu/myalu/_0813_ ), .A2(\myexu/myalu/_0765_ ), .A3(\myexu/myalu/_0797_ ), .ZN(\myexu/myalu/_0814_ ) );
BUF_X4 \myexu/myalu/_1797_ ( .A(\myexu/myalu/_0636_ ), .Z(\myexu/myalu/_0815_ ) );
AOI211_X2 \myexu/myalu/_1798_ ( .A(\myexu/myalu/_0798_ ), .B(\myexu/myalu/_0802_ ), .C1(\myexu/myalu/_0814_ ), .C2(\myexu/myalu/_0815_ ), .ZN(\myexu/myalu/_0816_ ) );
BUF_X4 \myexu/myalu/_1799_ ( .A(\myexu/myalu/_0726_ ), .Z(\myexu/myalu/_0817_ ) );
OAI21_X1 \myexu/myalu/_1800_ ( .A(\myexu/myalu/_0817_ ), .B1(fanout_net_11 ), .B2(\myexu/myalu/_1339_ ), .ZN(\myexu/myalu/_0818_ ) );
BUF_X4 \myexu/myalu/_1801_ ( .A(\myexu/myalu/_0721_ ), .Z(\myexu/myalu/_0819_ ) );
NAND2_X1 \myexu/myalu/_1802_ ( .A1(\myexu/myalu/_0496_ ), .A2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_0820_ ) );
BUF_X4 \myexu/myalu/_1803_ ( .A(\myexu/myalu/_0728_ ), .Z(\myexu/myalu/_0821_ ) );
BUF_X4 \myexu/myalu/_1804_ ( .A(\myexu/myalu/_0729_ ), .Z(\myexu/myalu/_0822_ ) );
AND2_X1 \myexu/myalu/_1805_ ( .A1(fanout_net_11 ), .A2(\myexu/myalu/_1339_ ), .ZN(\myexu/myalu/_0823_ ) );
NAND3_X1 \myexu/myalu/_1806_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0823_ ), .ZN(\myexu/myalu/_0824_ ) );
AND3_X1 \myexu/myalu/_1807_ ( .A1(\myexu/myalu/_0818_ ), .A2(\myexu/myalu/_0820_ ), .A3(\myexu/myalu/_0824_ ), .ZN(\myexu/myalu/_0825_ ) );
AND2_X4 \myexu/myalu/_1808_ ( .A1(\myexu/myalu/_0496_ ), .A2(\myexu/myalu/_0730_ ), .ZN(\myexu/myalu/_0826_ ) );
BUF_X2 \myexu/myalu/_1809_ ( .A(\myexu/myalu/_0723_ ), .Z(\myexu/myalu/_0827_ ) );
BUF_X4 \myexu/myalu/_1810_ ( .A(\myexu/myalu/_0827_ ), .Z(\myexu/myalu/_0828_ ) );
OAI21_X1 \myexu/myalu/_1811_ ( .A(\myexu/myalu/_0828_ ), .B1(\myexu/myalu/_0496_ ), .B2(\myexu/myalu/_0730_ ), .ZN(\myexu/myalu/_0829_ ) );
OAI211_X2 \myexu/myalu/_1812_ ( .A(\myexu/myalu/_0816_ ), .B(\myexu/myalu/_0825_ ), .C1(\myexu/myalu/_0826_ ), .C2(\myexu/myalu/_0829_ ), .ZN(\myexu/myalu/_1307_ ) );
BUF_X4 \myexu/myalu/_1813_ ( .A(\myexu/myalu/_0636_ ), .Z(\myexu/myalu/_0830_ ) );
INV_X1 \myexu/myalu/_1814_ ( .A(\myexu/myalu/_0812_ ), .ZN(\myexu/myalu/_0831_ ) );
NOR4_X1 \myexu/myalu/_1815_ ( .A1(\myexu/myalu/_0806_ ), .A2(\myexu/myalu/_0659_ ), .A3(\myexu/myalu/_0807_ ), .A4(\myexu/myalu/_0831_ ), .ZN(\myexu/myalu/_0832_ ) );
OAI21_X1 \myexu/myalu/_1816_ ( .A(\myexu/myalu/_0664_ ), .B1(\myexu/myalu/_0666_ ), .B2(\myexu/myalu/_0667_ ), .ZN(\myexu/myalu/_0833_ ) );
OAI21_X1 \myexu/myalu/_1817_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0643_ ), .B2(\myexu/myalu/_0644_ ), .ZN(\myexu/myalu/_0834_ ) );
AND3_X1 \myexu/myalu/_1818_ ( .A1(\myexu/myalu/_0833_ ), .A2(\myexu/myalu/_0834_ ), .A3(fanout_net_13 ), .ZN(\myexu/myalu/_0835_ ) );
NOR2_X1 \myexu/myalu/_1819_ ( .A1(\myexu/myalu/_0669_ ), .A2(\myexu/myalu/_0670_ ), .ZN(\myexu/myalu/_0836_ ) );
MUX2_X1 \myexu/myalu/_1820_ ( .A(\myexu/myalu/_0836_ ), .B(\myexu/myalu/_0663_ ), .S(\myexu/myalu/_0788_ ), .Z(\myexu/myalu/_0837_ ) );
AOI211_X4 \myexu/myalu/_1821_ ( .A(fanout_net_15 ), .B(\myexu/myalu/_0835_ ), .C1(\myexu/myalu/_0703_ ), .C2(\myexu/myalu/_0837_ ), .ZN(\myexu/myalu/_0838_ ) );
BUF_X4 \myexu/myalu/_1822_ ( .A(\myexu/myalu/_0788_ ), .Z(\myexu/myalu/_0839_ ) );
OAI21_X1 \myexu/myalu/_1823_ ( .A(\myexu/myalu/_0839_ ), .B1(\myexu/myalu/_0638_ ), .B2(\myexu/myalu/_0639_ ), .ZN(\myexu/myalu/_0840_ ) );
OAI21_X1 \myexu/myalu/_1824_ ( .A(fanout_net_11 ), .B1(\myexu/myalu/_0651_ ), .B2(\myexu/myalu/_0652_ ), .ZN(\myexu/myalu/_0841_ ) );
NAND2_X1 \myexu/myalu/_1825_ ( .A1(\myexu/myalu/_0840_ ), .A2(\myexu/myalu/_0841_ ), .ZN(\myexu/myalu/_0842_ ) );
BUF_X4 \myexu/myalu/_1826_ ( .A(\myexu/myalu/_0703_ ), .Z(\myexu/myalu/_0843_ ) );
NAND2_X1 \myexu/myalu/_1827_ ( .A1(\myexu/myalu/_0842_ ), .A2(\myexu/myalu/_0843_ ), .ZN(\myexu/myalu/_0844_ ) );
OR3_X1 \myexu/myalu/_1828_ ( .A1(\myexu/myalu/_0696_ ), .A2(\myexu/myalu/_0697_ ), .A3(\myexu/myalu/_0641_ ), .ZN(\myexu/myalu/_0845_ ) );
OR3_X1 \myexu/myalu/_1829_ ( .A1(\myexu/myalu/_0648_ ), .A2(\myexu/myalu/_0649_ ), .A3(fanout_net_11 ), .ZN(\myexu/myalu/_0846_ ) );
NAND3_X1 \myexu/myalu/_1830_ ( .A1(\myexu/myalu/_0845_ ), .A2(\myexu/myalu/_0846_ ), .A3(fanout_net_13 ), .ZN(\myexu/myalu/_0847_ ) );
NAND2_X1 \myexu/myalu/_1831_ ( .A1(\myexu/myalu/_0844_ ), .A2(\myexu/myalu/_0847_ ), .ZN(\myexu/myalu/_0848_ ) );
AOI211_X4 \myexu/myalu/_1832_ ( .A(fanout_net_17 ), .B(\myexu/myalu/_0838_ ), .C1(fanout_net_15 ), .C2(\myexu/myalu/_0848_ ), .ZN(\myexu/myalu/_0849_ ) );
OAI21_X1 \myexu/myalu/_1833_ ( .A(\myexu/myalu/_0664_ ), .B1(\myexu/myalu/_0699_ ), .B2(\myexu/myalu/_0700_ ), .ZN(\myexu/myalu/_0850_ ) );
OAI21_X1 \myexu/myalu/_1834_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0705_ ), .B2(\myexu/myalu/_0706_ ), .ZN(\myexu/myalu/_0851_ ) );
NAND2_X1 \myexu/myalu/_1835_ ( .A1(\myexu/myalu/_0850_ ), .A2(\myexu/myalu/_0851_ ), .ZN(\myexu/myalu/_0852_ ) );
NAND2_X1 \myexu/myalu/_1836_ ( .A1(\myexu/myalu/_0852_ ), .A2(\myexu/myalu/_0773_ ), .ZN(\myexu/myalu/_0853_ ) );
OR3_X1 \myexu/myalu/_1837_ ( .A1(\myexu/myalu/_0683_ ), .A2(\myexu/myalu/_0684_ ), .A3(\myexu/myalu/_0641_ ), .ZN(\myexu/myalu/_0854_ ) );
INV_X1 \myexu/myalu/_1838_ ( .A(\myexu/myalu/_0709_ ), .ZN(\myexu/myalu/_0855_ ) );
OAI211_X2 \myexu/myalu/_1839_ ( .A(\myexu/myalu/_0855_ ), .B(\myexu/myalu/_0788_ ), .C1(fanout_net_10 ), .C2(\myexu/myalu/_0545_ ), .ZN(\myexu/myalu/_0856_ ) );
NAND3_X1 \myexu/myalu/_1840_ ( .A1(\myexu/myalu/_0854_ ), .A2(\myexu/myalu/_0856_ ), .A3(fanout_net_13 ), .ZN(\myexu/myalu/_0857_ ) );
NAND2_X1 \myexu/myalu/_1841_ ( .A1(\myexu/myalu/_0853_ ), .A2(\myexu/myalu/_0857_ ), .ZN(\myexu/myalu/_0858_ ) );
OAI21_X1 \myexu/myalu/_1842_ ( .A(\myexu/myalu/_0641_ ), .B1(\myexu/myalu/_0679_ ), .B2(\myexu/myalu/_0680_ ), .ZN(\myexu/myalu/_0859_ ) );
OAI21_X1 \myexu/myalu/_1843_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0689_ ), .B2(\myexu/myalu/_0690_ ), .ZN(\myexu/myalu/_0860_ ) );
NAND2_X1 \myexu/myalu/_1844_ ( .A1(\myexu/myalu/_0859_ ), .A2(\myexu/myalu/_0860_ ), .ZN(\myexu/myalu/_0861_ ) );
AND2_X1 \myexu/myalu/_1845_ ( .A1(\myexu/myalu/_0687_ ), .A2(\myexu/myalu/_0664_ ), .ZN(\myexu/myalu/_0862_ ) );
MUX2_X1 \myexu/myalu/_1846_ ( .A(\myexu/myalu/_0861_ ), .B(\myexu/myalu/_0862_ ), .S(fanout_net_13 ), .Z(\myexu/myalu/_0863_ ) );
MUX2_X1 \myexu/myalu/_1847_ ( .A(\myexu/myalu/_0858_ ), .B(\myexu/myalu/_0863_ ), .S(fanout_net_15 ), .Z(\myexu/myalu/_0864_ ) );
BUF_X4 \myexu/myalu/_1848_ ( .A(\myexu/myalu/_0588_ ), .Z(\myexu/myalu/_0865_ ) );
BUF_X4 \myexu/myalu/_1849_ ( .A(\myexu/myalu/_0865_ ), .Z(\myexu/myalu/_0866_ ) );
BUF_X4 \myexu/myalu/_1850_ ( .A(\myexu/myalu/_0866_ ), .Z(\myexu/myalu/_0867_ ) );
NOR2_X1 \myexu/myalu/_1851_ ( .A1(\myexu/myalu/_0864_ ), .A2(\myexu/myalu/_0867_ ), .ZN(\myexu/myalu/_0868_ ) );
NOR2_X1 \myexu/myalu/_1852_ ( .A1(\myexu/myalu/_0849_ ), .A2(\myexu/myalu/_0868_ ), .ZN(\myexu/myalu/_0869_ ) );
OAI21_X1 \myexu/myalu/_1853_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_0832_ ), .B2(\myexu/myalu/_0869_ ), .ZN(\myexu/myalu/_0870_ ) );
OR3_X1 \myexu/myalu/_1854_ ( .A1(\myexu/myalu/_0849_ ), .A2(\myexu/myalu/_0734_ ), .A3(\myexu/myalu/_0868_ ), .ZN(\myexu/myalu/_0871_ ) );
INV_X1 \myexu/myalu/_1855_ ( .A(\myexu/myalu/_0726_ ), .ZN(\myexu/myalu/_0872_ ) );
BUF_X4 \myexu/myalu/_1856_ ( .A(\myexu/myalu/_0843_ ), .Z(\myexu/myalu/_0873_ ) );
AOI21_X1 \myexu/myalu/_1857_ ( .A(\myexu/myalu/_0872_ ), .B1(\myexu/myalu/_0873_ ), .B2(\myexu/myalu/_0502_ ), .ZN(\myexu/myalu/_0874_ ) );
BUF_X4 \myexu/myalu/_1858_ ( .A(\myexu/myalu/_0721_ ), .Z(\myexu/myalu/_0875_ ) );
NAND3_X1 \myexu/myalu/_1859_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_1328_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0876_ ) );
AND2_X1 \myexu/myalu/_1860_ ( .A1(\myexu/myalu/_1360_ ), .A2(\myexu/myalu/_1339_ ), .ZN(\myexu/myalu/_0877_ ) );
NOR2_X1 \myexu/myalu/_1861_ ( .A1(\myexu/myalu/_0661_ ), .A2(\myexu/myalu/_0877_ ), .ZN(\myexu/myalu/_0878_ ) );
OAI21_X1 \myexu/myalu/_1862_ ( .A(\myexu/myalu/_0876_ ), .B1(\myexu/myalu/_0878_ ), .B2(fanout_net_12 ), .ZN(\myexu/myalu/_0879_ ) );
BUF_X2 \myexu/myalu/_1863_ ( .A(\myexu/myalu/_0646_ ), .Z(\myexu/myalu/_0880_ ) );
AND2_X1 \myexu/myalu/_1864_ ( .A1(\myexu/myalu/_0879_ ), .A2(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_0881_ ) );
BUF_X4 \myexu/myalu/_1865_ ( .A(\myexu/myalu/_0506_ ), .Z(\myexu/myalu/_0882_ ) );
BUF_X4 \myexu/myalu/_1866_ ( .A(\myexu/myalu/_0882_ ), .Z(\myexu/myalu/_0883_ ) );
AND2_X1 \myexu/myalu/_1867_ ( .A1(\myexu/myalu/_0881_ ), .A2(\myexu/myalu/_0883_ ), .ZN(\myexu/myalu/_0884_ ) );
BUF_X4 \myexu/myalu/_1868_ ( .A(\myexu/myalu/_0718_ ), .Z(\myexu/myalu/_0885_ ) );
BUF_X4 \myexu/myalu/_1869_ ( .A(\myexu/myalu/_0885_ ), .Z(\myexu/myalu/_0886_ ) );
AOI221_X4 \myexu/myalu/_1870_ ( .A(\myexu/myalu/_0874_ ), .B1(\myexu/myalu/_0494_ ), .B2(\myexu/myalu/_0875_ ), .C1(\myexu/myalu/_0884_ ), .C2(\myexu/myalu/_0886_ ), .ZN(\myexu/myalu/_0887_ ) );
NOR2_X1 \myexu/myalu/_1871_ ( .A1(\myexu/myalu/_0826_ ), .A2(\myexu/myalu/_0823_ ), .ZN(\myexu/myalu/_0888_ ) );
AOI21_X1 \myexu/myalu/_1872_ ( .A(\myexu/myalu/_0724_ ), .B1(\myexu/myalu/_0888_ ), .B2(\myexu/myalu/_0495_ ), .ZN(\myexu/myalu/_0889_ ) );
OAI21_X1 \myexu/myalu/_1873_ ( .A(\myexu/myalu/_0889_ ), .B1(\myexu/myalu/_0495_ ), .B2(\myexu/myalu/_0888_ ), .ZN(\myexu/myalu/_0890_ ) );
AND2_X1 \myexu/myalu/_1874_ ( .A1(fanout_net_13 ), .A2(\myexu/myalu/_1350_ ), .ZN(\myexu/myalu/_0891_ ) );
NAND3_X1 \myexu/myalu/_1875_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0891_ ), .ZN(\myexu/myalu/_0892_ ) );
AND2_X1 \myexu/myalu/_1876_ ( .A1(\myexu/myalu/_0890_ ), .A2(\myexu/myalu/_0892_ ), .ZN(\myexu/myalu/_0893_ ) );
NAND4_X1 \myexu/myalu/_1877_ ( .A1(\myexu/myalu/_0870_ ), .A2(\myexu/myalu/_0871_ ), .A3(\myexu/myalu/_0887_ ), .A4(\myexu/myalu/_0893_ ), .ZN(\myexu/myalu/_1318_ ) );
NOR3_X1 \myexu/myalu/_1878_ ( .A1(\myexu/myalu/_0806_ ), .A2(\myexu/myalu/_0807_ ), .A3(\myexu/myalu/_0831_ ), .ZN(\myexu/myalu/_0894_ ) );
OR3_X1 \myexu/myalu/_1879_ ( .A1(\myexu/myalu/_0756_ ), .A2(\myexu/myalu/_0664_ ), .A3(\myexu/myalu/_0757_ ), .ZN(\myexu/myalu/_0895_ ) );
OR3_X1 \myexu/myalu/_1880_ ( .A1(\myexu/myalu/_0743_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0744_ ), .ZN(\myexu/myalu/_0896_ ) );
NAND3_X1 \myexu/myalu/_1881_ ( .A1(\myexu/myalu/_0895_ ), .A2(\myexu/myalu/_0896_ ), .A3(fanout_net_13 ), .ZN(\myexu/myalu/_0897_ ) );
OR3_X1 \myexu/myalu/_1882_ ( .A1(\myexu/myalu/_0735_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0736_ ), .ZN(\myexu/myalu/_0898_ ) );
OR3_X1 \myexu/myalu/_1883_ ( .A1(\myexu/myalu/_0746_ ), .A2(\myexu/myalu/_0747_ ), .A3(\myexu/myalu/_0641_ ), .ZN(\myexu/myalu/_0899_ ) );
NAND3_X1 \myexu/myalu/_1884_ ( .A1(\myexu/myalu/_0898_ ), .A2(\myexu/myalu/_0773_ ), .A3(\myexu/myalu/_0899_ ), .ZN(\myexu/myalu/_0900_ ) );
AND3_X1 \myexu/myalu/_1885_ ( .A1(\myexu/myalu/_0897_ ), .A2(\myexu/myalu/_0900_ ), .A3(\myexu/myalu/_0506_ ), .ZN(\myexu/myalu/_0901_ ) );
NAND2_X1 \myexu/myalu/_1886_ ( .A1(\myexu/myalu/_0754_ ), .A2(fanout_net_12 ), .ZN(\myexu/myalu/_0902_ ) );
OR3_X1 \myexu/myalu/_1887_ ( .A1(\myexu/myalu/_0759_ ), .A2(\myexu/myalu/_0760_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0903_ ) );
NAND3_X1 \myexu/myalu/_1888_ ( .A1(\myexu/myalu/_0902_ ), .A2(\myexu/myalu/_0903_ ), .A3(\myexu/myalu/_0773_ ), .ZN(\myexu/myalu/_0904_ ) );
BUF_X2 \myexu/myalu/_1889_ ( .A(\myexu/myalu/_0788_ ), .Z(\myexu/myalu/_0905_ ) );
NAND4_X1 \myexu/myalu/_1890_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_0905_ ), .A3(fanout_net_13 ), .A4(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_0906_ ) );
AND2_X1 \myexu/myalu/_1891_ ( .A1(\myexu/myalu/_0904_ ), .A2(\myexu/myalu/_0906_ ), .ZN(\myexu/myalu/_0907_ ) );
AOI21_X1 \myexu/myalu/_1892_ ( .A(\myexu/myalu/_0901_ ), .B1(fanout_net_15 ), .B2(\myexu/myalu/_0907_ ), .ZN(\myexu/myalu/_0908_ ) );
NAND2_X1 \myexu/myalu/_1893_ ( .A1(\myexu/myalu/_0908_ ), .A2(fanout_net_17 ), .ZN(\myexu/myalu/_0909_ ) );
BUF_X4 \myexu/myalu/_1894_ ( .A(\myexu/myalu/_0865_ ), .Z(\myexu/myalu/_0910_ ) );
BUF_X4 \myexu/myalu/_1895_ ( .A(\myexu/myalu/_0910_ ), .Z(\myexu/myalu/_0911_ ) );
OR3_X1 \myexu/myalu/_1896_ ( .A1(\myexu/myalu/_0766_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0767_ ), .ZN(\myexu/myalu/_0912_ ) );
OR3_X1 \myexu/myalu/_1897_ ( .A1(\myexu/myalu/_0778_ ), .A2(\myexu/myalu/_0779_ ), .A3(\myexu/myalu/_0664_ ), .ZN(\myexu/myalu/_0913_ ) );
NAND3_X1 \myexu/myalu/_1898_ ( .A1(\myexu/myalu/_0912_ ), .A2(\myexu/myalu/_0880_ ), .A3(\myexu/myalu/_0913_ ), .ZN(\myexu/myalu/_0914_ ) );
OR3_X1 \myexu/myalu/_1899_ ( .A1(\myexu/myalu/_0775_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0776_ ), .ZN(\myexu/myalu/_0915_ ) );
OR3_X1 \myexu/myalu/_1900_ ( .A1(\myexu/myalu/_0738_ ), .A2(\myexu/myalu/_0739_ ), .A3(\myexu/myalu/_0788_ ), .ZN(\myexu/myalu/_0916_ ) );
NAND3_X1 \myexu/myalu/_1901_ ( .A1(\myexu/myalu/_0915_ ), .A2(fanout_net_13 ), .A3(\myexu/myalu/_0916_ ), .ZN(\myexu/myalu/_0917_ ) );
NAND3_X1 \myexu/myalu/_1902_ ( .A1(\myexu/myalu/_0914_ ), .A2(\myexu/myalu/_0917_ ), .A3(fanout_net_15 ), .ZN(\myexu/myalu/_0918_ ) );
OAI21_X1 \myexu/myalu/_1903_ ( .A(\myexu/myalu/_0905_ ), .B1(\myexu/myalu/_0792_ ), .B2(\myexu/myalu/_0793_ ), .ZN(\myexu/myalu/_0919_ ) );
OAI21_X1 \myexu/myalu/_1904_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0769_ ), .B2(\myexu/myalu/_0770_ ), .ZN(\myexu/myalu/_0920_ ) );
NAND2_X1 \myexu/myalu/_1905_ ( .A1(\myexu/myalu/_0919_ ), .A2(\myexu/myalu/_0920_ ), .ZN(\myexu/myalu/_0921_ ) );
NOR3_X1 \myexu/myalu/_1906_ ( .A1(\myexu/myalu/_0789_ ), .A2(\myexu/myalu/_0839_ ), .A3(\myexu/myalu/_0790_ ), .ZN(\myexu/myalu/_0922_ ) );
NOR3_X1 \myexu/myalu/_1907_ ( .A1(\myexu/myalu/_0783_ ), .A2(\myexu/myalu/_0784_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0923_ ) );
NOR2_X1 \myexu/myalu/_1908_ ( .A1(\myexu/myalu/_0922_ ), .A2(\myexu/myalu/_0923_ ), .ZN(\myexu/myalu/_0924_ ) );
MUX2_X1 \myexu/myalu/_1909_ ( .A(\myexu/myalu/_0921_ ), .B(\myexu/myalu/_0924_ ), .S(\myexu/myalu/_0873_ ), .Z(\myexu/myalu/_0925_ ) );
OAI211_X2 \myexu/myalu/_1910_ ( .A(\myexu/myalu/_0911_ ), .B(\myexu/myalu/_0918_ ), .C1(\myexu/myalu/_0925_ ), .C2(fanout_net_15 ), .ZN(\myexu/myalu/_0926_ ) );
NAND2_X1 \myexu/myalu/_1911_ ( .A1(\myexu/myalu/_0909_ ), .A2(\myexu/myalu/_0926_ ), .ZN(\myexu/myalu/_0927_ ) );
OAI21_X1 \myexu/myalu/_1912_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_0894_ ), .B2(\myexu/myalu/_0927_ ), .ZN(\myexu/myalu/_0928_ ) );
BUF_X2 \myexu/myalu/_1913_ ( .A(\myexu/myalu/_0677_ ), .Z(\myexu/myalu/_0929_ ) );
BUF_X2 \myexu/myalu/_1914_ ( .A(\myexu/myalu/_0929_ ), .Z(\myexu/myalu/_0930_ ) );
NAND2_X1 \myexu/myalu/_1915_ ( .A1(\myexu/myalu/_0927_ ), .A2(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0931_ ) );
BUF_X4 \myexu/myalu/_1916_ ( .A(\myexu/myalu/_0724_ ), .Z(\myexu/myalu/_0932_ ) );
NOR2_X1 \myexu/myalu/_1917_ ( .A1(\myexu/myalu/_0888_ ), .A2(\myexu/myalu/_0495_ ), .ZN(\myexu/myalu/_0933_ ) );
NOR2_X1 \myexu/myalu/_1918_ ( .A1(\myexu/myalu/_0933_ ), .A2(\myexu/myalu/_0891_ ), .ZN(\myexu/myalu/_0934_ ) );
AOI21_X1 \myexu/myalu/_1919_ ( .A(\myexu/myalu/_0932_ ), .B1(\myexu/myalu/_0934_ ), .B2(\myexu/myalu/_0493_ ), .ZN(\myexu/myalu/_0935_ ) );
OAI21_X1 \myexu/myalu/_1920_ ( .A(\myexu/myalu/_0935_ ), .B1(\myexu/myalu/_0493_ ), .B2(\myexu/myalu/_0934_ ), .ZN(\myexu/myalu/_0936_ ) );
OAI21_X1 \myexu/myalu/_1921_ ( .A(\myexu/myalu/_0817_ ), .B1(fanout_net_15 ), .B2(\myexu/myalu/_1353_ ), .ZN(\myexu/myalu/_0937_ ) );
AND2_X1 \myexu/myalu/_1922_ ( .A1(\myexu/myalu/_1360_ ), .A2(\myexu/myalu/_1350_ ), .ZN(\myexu/myalu/_0938_ ) );
NOR2_X1 \myexu/myalu/_1923_ ( .A1(\myexu/myalu/_0783_ ), .A2(\myexu/myalu/_0938_ ), .ZN(\myexu/myalu/_0939_ ) );
MUX2_X1 \myexu/myalu/_1924_ ( .A(\myexu/myalu/_0799_ ), .B(\myexu/myalu/_0939_ ), .S(\myexu/myalu/_0695_ ), .Z(\myexu/myalu/_0940_ ) );
OR2_X1 \myexu/myalu/_1925_ ( .A1(\myexu/myalu/_0940_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0941_ ) );
INV_X1 \myexu/myalu/_1926_ ( .A(\myexu/myalu/_0718_ ), .ZN(\myexu/myalu/_0942_ ) );
OR3_X1 \myexu/myalu/_1927_ ( .A1(\myexu/myalu/_0941_ ), .A2(fanout_net_15 ), .A3(\myexu/myalu/_0942_ ), .ZN(\myexu/myalu/_0943_ ) );
BUF_X2 \myexu/myalu/_1928_ ( .A(\myexu/myalu/_0728_ ), .Z(\myexu/myalu/_0944_ ) );
BUF_X4 \myexu/myalu/_1929_ ( .A(\myexu/myalu/_0729_ ), .Z(\myexu/myalu/_0945_ ) );
AND2_X1 \myexu/myalu/_1930_ ( .A1(fanout_net_15 ), .A2(\myexu/myalu/_1353_ ), .ZN(\myexu/myalu/_0946_ ) );
NAND3_X1 \myexu/myalu/_1931_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0946_ ), .ZN(\myexu/myalu/_0947_ ) );
OR2_X1 \myexu/myalu/_1932_ ( .A1(\myexu/myalu/_0722_ ), .A2(\myexu/myalu/_0493_ ), .ZN(\myexu/myalu/_0948_ ) );
AND4_X1 \myexu/myalu/_1933_ ( .A1(\myexu/myalu/_0937_ ), .A2(\myexu/myalu/_0943_ ), .A3(\myexu/myalu/_0947_ ), .A4(\myexu/myalu/_0948_ ), .ZN(\myexu/myalu/_0949_ ) );
NAND4_X1 \myexu/myalu/_1934_ ( .A1(\myexu/myalu/_0928_ ), .A2(\myexu/myalu/_0931_ ), .A3(\myexu/myalu/_0936_ ), .A4(\myexu/myalu/_0949_ ), .ZN(\myexu/myalu/_1321_ ) );
INV_X2 \myexu/myalu/_1935_ ( .A(\myexu/myalu/_0636_ ), .ZN(\myexu/myalu/_0950_ ) );
NAND4_X1 \myexu/myalu/_1936_ ( .A1(\myexu/myalu/_0634_ ), .A2(\myexu/myalu/_0803_ ), .A3(\myexu/myalu/_0805_ ), .A4(\myexu/myalu/_0812_ ), .ZN(\myexu/myalu/_0951_ ) );
AOI21_X1 \myexu/myalu/_1937_ ( .A(\myexu/myalu/_0646_ ), .B1(\myexu/myalu/_0681_ ), .B2(\myexu/myalu/_0685_ ), .ZN(\myexu/myalu/_0952_ ) );
AND3_X1 \myexu/myalu/_1938_ ( .A1(\myexu/myalu/_0707_ ), .A2(\myexu/myalu/_0710_ ), .A3(\myexu/myalu/_0646_ ), .ZN(\myexu/myalu/_0953_ ) );
OR3_X1 \myexu/myalu/_1939_ ( .A1(\myexu/myalu/_0952_ ), .A2(\myexu/myalu/_0953_ ), .A3(fanout_net_15 ), .ZN(\myexu/myalu/_0954_ ) );
NAND4_X1 \myexu/myalu/_1940_ ( .A1(\myexu/myalu/_0688_ ), .A2(fanout_net_15 ), .A3(\myexu/myalu/_0703_ ), .A4(\myexu/myalu/_0691_ ), .ZN(\myexu/myalu/_0955_ ) );
NAND2_X1 \myexu/myalu/_1941_ ( .A1(\myexu/myalu/_0954_ ), .A2(\myexu/myalu/_0955_ ), .ZN(\myexu/myalu/_0956_ ) );
NAND2_X1 \myexu/myalu/_1942_ ( .A1(\myexu/myalu/_0956_ ), .A2(fanout_net_17 ), .ZN(\myexu/myalu/_0957_ ) );
NAND2_X1 \myexu/myalu/_1943_ ( .A1(\myexu/myalu/_0702_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0958_ ) );
NAND3_X1 \myexu/myalu/_1944_ ( .A1(\myexu/myalu/_0650_ ), .A2(\myexu/myalu/_0653_ ), .A3(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_0959_ ) );
NAND3_X1 \myexu/myalu/_1945_ ( .A1(\myexu/myalu/_0958_ ), .A2(\myexu/myalu/_0959_ ), .A3(fanout_net_15 ), .ZN(\myexu/myalu/_0960_ ) );
AND2_X1 \myexu/myalu/_1946_ ( .A1(\myexu/myalu/_0642_ ), .A2(\myexu/myalu/_0645_ ), .ZN(\myexu/myalu/_0961_ ) );
MUX2_X1 \myexu/myalu/_1947_ ( .A(\myexu/myalu/_0672_ ), .B(\myexu/myalu/_0961_ ), .S(fanout_net_13 ), .Z(\myexu/myalu/_0962_ ) );
OAI211_X2 \myexu/myalu/_1948_ ( .A(\myexu/myalu/_0866_ ), .B(\myexu/myalu/_0960_ ), .C1(\myexu/myalu/_0962_ ), .C2(fanout_net_15 ), .ZN(\myexu/myalu/_0963_ ) );
AND2_X1 \myexu/myalu/_1949_ ( .A1(\myexu/myalu/_0957_ ), .A2(\myexu/myalu/_0963_ ), .ZN(\myexu/myalu/_0964_ ) );
AOI21_X1 \myexu/myalu/_1950_ ( .A(\myexu/myalu/_0950_ ), .B1(\myexu/myalu/_0951_ ), .B2(\myexu/myalu/_0964_ ), .ZN(\myexu/myalu/_0965_ ) );
AOI21_X1 \myexu/myalu/_1951_ ( .A(\myexu/myalu/_0734_ ), .B1(\myexu/myalu/_0957_ ), .B2(\myexu/myalu/_0963_ ), .ZN(\myexu/myalu/_0966_ ) );
NOR3_X2 \myexu/myalu/_1952_ ( .A1(\myexu/myalu/_0888_ ), .A2(\myexu/myalu/_0493_ ), .A3(\myexu/myalu/_0495_ ), .ZN(\myexu/myalu/_0967_ ) );
NOR3_X1 \myexu/myalu/_1953_ ( .A1(\myexu/myalu/_0493_ ), .A2(\myexu/myalu/_0585_ ), .A3(\myexu/myalu/_0502_ ), .ZN(\myexu/myalu/_0968_ ) );
OR2_X1 \myexu/myalu/_1954_ ( .A1(\myexu/myalu/_0968_ ), .A2(\myexu/myalu/_0946_ ), .ZN(\myexu/myalu/_0969_ ) );
NOR2_X1 \myexu/myalu/_1955_ ( .A1(\myexu/myalu/_0967_ ), .A2(\myexu/myalu/_0969_ ), .ZN(\myexu/myalu/_0970_ ) );
INV_X1 \myexu/myalu/_1956_ ( .A(\myexu/myalu/_0970_ ), .ZN(\myexu/myalu/_0971_ ) );
AND2_X1 \myexu/myalu/_1957_ ( .A1(\myexu/myalu/_0971_ ), .A2(\myexu/myalu/_0491_ ), .ZN(\myexu/myalu/_0972_ ) );
OAI21_X1 \myexu/myalu/_1958_ ( .A(\myexu/myalu/_0827_ ), .B1(\myexu/myalu/_0971_ ), .B2(\myexu/myalu/_0491_ ), .ZN(\myexu/myalu/_0973_ ) );
NOR2_X1 \myexu/myalu/_1959_ ( .A1(\myexu/myalu/_0972_ ), .A2(\myexu/myalu/_0973_ ), .ZN(\myexu/myalu/_0974_ ) );
NAND4_X1 \myexu/myalu/_1960_ ( .A1(\myexu/myalu/_0658_ ), .A2(\myexu/myalu/_0839_ ), .A3(\myexu/myalu/_1328_ ), .A4(fanout_net_13 ), .ZN(\myexu/myalu/_0975_ ) );
OAI21_X1 \myexu/myalu/_1961_ ( .A(\myexu/myalu/_0839_ ), .B1(\myexu/myalu/_0669_ ), .B2(\myexu/myalu/_0662_ ), .ZN(\myexu/myalu/_0976_ ) );
OAI21_X1 \myexu/myalu/_1962_ ( .A(\myexu/myalu/_0976_ ), .B1(\myexu/myalu/_0878_ ), .B2(\myexu/myalu/_0839_ ), .ZN(\myexu/myalu/_0977_ ) );
INV_X1 \myexu/myalu/_1963_ ( .A(\myexu/myalu/_0977_ ), .ZN(\myexu/myalu/_0978_ ) );
OAI21_X1 \myexu/myalu/_1964_ ( .A(\myexu/myalu/_0975_ ), .B1(\myexu/myalu/_0978_ ), .B2(fanout_net_13 ), .ZN(\myexu/myalu/_0979_ ) );
BUF_X4 \myexu/myalu/_1965_ ( .A(\myexu/myalu/_0883_ ), .Z(\myexu/myalu/_0980_ ) );
NAND3_X1 \myexu/myalu/_1966_ ( .A1(\myexu/myalu/_0979_ ), .A2(\myexu/myalu/_0980_ ), .A3(\myexu/myalu/_0885_ ), .ZN(\myexu/myalu/_0981_ ) );
NAND2_X1 \myexu/myalu/_1967_ ( .A1(\myexu/myalu/_0491_ ), .A2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0982_ ) );
BUF_X4 \myexu/myalu/_1968_ ( .A(\myexu/myalu/_0729_ ), .Z(\myexu/myalu/_0983_ ) );
AND2_X1 \myexu/myalu/_1969_ ( .A1(fanout_net_17 ), .A2(\myexu/myalu/_1354_ ), .ZN(\myexu/myalu/_0984_ ) );
NAND3_X1 \myexu/myalu/_1970_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0984_ ), .ZN(\myexu/myalu/_0985_ ) );
OAI21_X1 \myexu/myalu/_1971_ ( .A(\myexu/myalu/_0817_ ), .B1(fanout_net_17 ), .B2(\myexu/myalu/_1354_ ), .ZN(\myexu/myalu/_0986_ ) );
NAND4_X1 \myexu/myalu/_1972_ ( .A1(\myexu/myalu/_0981_ ), .A2(\myexu/myalu/_0982_ ), .A3(\myexu/myalu/_0985_ ), .A4(\myexu/myalu/_0986_ ), .ZN(\myexu/myalu/_0987_ ) );
OR4_X1 \myexu/myalu/_1973_ ( .A1(\myexu/myalu/_0965_ ), .A2(\myexu/myalu/_0966_ ), .A3(\myexu/myalu/_0974_ ), .A4(\myexu/myalu/_0987_ ), .ZN(\myexu/myalu/_1322_ ) );
AND2_X1 \myexu/myalu/_1974_ ( .A1(\myexu/myalu/_0755_ ), .A2(\myexu/myalu/_0773_ ), .ZN(\myexu/myalu/_0988_ ) );
NAND2_X1 \myexu/myalu/_1975_ ( .A1(\myexu/myalu/_0749_ ), .A2(\myexu/myalu/_0646_ ), .ZN(\myexu/myalu/_0989_ ) );
NAND2_X1 \myexu/myalu/_1976_ ( .A1(\myexu/myalu/_0762_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_0990_ ) );
NAND2_X1 \myexu/myalu/_1977_ ( .A1(\myexu/myalu/_0989_ ), .A2(\myexu/myalu/_0990_ ), .ZN(\myexu/myalu/_0991_ ) );
MUX2_X1 \myexu/myalu/_1978_ ( .A(\myexu/myalu/_0988_ ), .B(\myexu/myalu/_0991_ ), .S(\myexu/myalu/_0506_ ), .Z(\myexu/myalu/_0992_ ) );
OR2_X1 \myexu/myalu/_1979_ ( .A1(\myexu/myalu/_0992_ ), .A2(\myexu/myalu/_0866_ ), .ZN(\myexu/myalu/_0993_ ) );
NAND3_X1 \myexu/myalu/_1980_ ( .A1(\myexu/myalu/_0791_ ), .A2(\myexu/myalu/_0843_ ), .A3(\myexu/myalu/_0794_ ), .ZN(\myexu/myalu/_0994_ ) );
BUF_X4 \myexu/myalu/_1981_ ( .A(\myexu/myalu/_0506_ ), .Z(\myexu/myalu/_0995_ ) );
BUF_X4 \myexu/myalu/_1982_ ( .A(\myexu/myalu/_0703_ ), .Z(\myexu/myalu/_0996_ ) );
OAI211_X2 \myexu/myalu/_1983_ ( .A(\myexu/myalu/_0994_ ), .B(\myexu/myalu/_0995_ ), .C1(\myexu/myalu/_0772_ ), .C2(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_0997_ ) );
AND3_X1 \myexu/myalu/_1984_ ( .A1(\myexu/myalu/_0777_ ), .A2(\myexu/myalu/_0646_ ), .A3(\myexu/myalu/_0780_ ), .ZN(\myexu/myalu/_0998_ ) );
AOI21_X1 \myexu/myalu/_1985_ ( .A(\myexu/myalu/_0998_ ), .B1(fanout_net_13 ), .B2(\myexu/myalu/_0741_ ), .ZN(\myexu/myalu/_0999_ ) );
BUF_X4 \myexu/myalu/_1986_ ( .A(\myexu/myalu/_0995_ ), .Z(\myexu/myalu/_1000_ ) );
OAI211_X2 \myexu/myalu/_1987_ ( .A(\myexu/myalu/_0910_ ), .B(\myexu/myalu/_0997_ ), .C1(\myexu/myalu/_0999_ ), .C2(\myexu/myalu/_1000_ ), .ZN(\myexu/myalu/_1001_ ) );
AND3_X1 \myexu/myalu/_1988_ ( .A1(\myexu/myalu/_0993_ ), .A2(\myexu/myalu/_0930_ ), .A3(\myexu/myalu/_1001_ ), .ZN(\myexu/myalu/_1002_ ) );
OR2_X2 \myexu/myalu/_1989_ ( .A1(\myexu/myalu/_0809_ ), .A2(fanout_net_13 ), .ZN(\myexu/myalu/_1003_ ) );
NAND4_X1 \myexu/myalu/_1990_ ( .A1(\myexu/myalu/_0634_ ), .A2(\myexu/myalu/_0803_ ), .A3(\myexu/myalu/_0812_ ), .A4(\myexu/myalu/_1003_ ), .ZN(\myexu/myalu/_1004_ ) );
NAND2_X1 \myexu/myalu/_1991_ ( .A1(\myexu/myalu/_0993_ ), .A2(\myexu/myalu/_1001_ ), .ZN(\myexu/myalu/_1005_ ) );
AOI21_X1 \myexu/myalu/_1992_ ( .A(\myexu/myalu/_0950_ ), .B1(\myexu/myalu/_1004_ ), .B2(\myexu/myalu/_1005_ ), .ZN(\myexu/myalu/_1006_ ) );
OR3_X1 \myexu/myalu/_1993_ ( .A1(\myexu/myalu/_0972_ ), .A2(\myexu/myalu/_0482_ ), .A3(\myexu/myalu/_0984_ ), .ZN(\myexu/myalu/_1007_ ) );
OAI21_X1 \myexu/myalu/_1994_ ( .A(\myexu/myalu/_0482_ ), .B1(\myexu/myalu/_0972_ ), .B2(\myexu/myalu/_0984_ ), .ZN(\myexu/myalu/_1008_ ) );
AND3_X1 \myexu/myalu/_1995_ ( .A1(\myexu/myalu/_1007_ ), .A2(\myexu/myalu/_0827_ ), .A3(\myexu/myalu/_1008_ ), .ZN(\myexu/myalu/_1009_ ) );
NOR2_X1 \myexu/myalu/_1996_ ( .A1(\myexu/myalu/_0799_ ), .A2(fanout_net_12 ), .ZN(\myexu/myalu/_1010_ ) );
OR3_X1 \myexu/myalu/_1997_ ( .A1(\myexu/myalu/_0789_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0784_ ), .ZN(\myexu/myalu/_1011_ ) );
OR3_X1 \myexu/myalu/_1998_ ( .A1(\myexu/myalu/_0783_ ), .A2(\myexu/myalu/_0938_ ), .A3(\myexu/myalu/_0664_ ), .ZN(\myexu/myalu/_1012_ ) );
AND2_X1 \myexu/myalu/_1999_ ( .A1(\myexu/myalu/_1011_ ), .A2(\myexu/myalu/_1012_ ), .ZN(\myexu/myalu/_1013_ ) );
MUX2_X1 \myexu/myalu/_2000_ ( .A(\myexu/myalu/_1010_ ), .B(\myexu/myalu/_1013_ ), .S(\myexu/myalu/_0703_ ), .Z(\myexu/myalu/_1014_ ) );
NAND3_X1 \myexu/myalu/_2001_ ( .A1(\myexu/myalu/_1014_ ), .A2(\myexu/myalu/_0980_ ), .A3(\myexu/myalu/_0885_ ), .ZN(\myexu/myalu/_1015_ ) );
NAND2_X1 \myexu/myalu/_2002_ ( .A1(\myexu/myalu/_0482_ ), .A2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_1016_ ) );
AND2_X1 \myexu/myalu/_2003_ ( .A1(\myexu/myalu/_1387_ ), .A2(\myexu/myalu/_1355_ ), .ZN(\myexu/myalu/_1017_ ) );
NAND3_X1 \myexu/myalu/_2004_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0729_ ), .A3(\myexu/myalu/_1017_ ), .ZN(\myexu/myalu/_1018_ ) );
OAI21_X1 \myexu/myalu/_2005_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1387_ ), .B2(\myexu/myalu/_1355_ ), .ZN(\myexu/myalu/_1019_ ) );
NAND4_X1 \myexu/myalu/_2006_ ( .A1(\myexu/myalu/_1015_ ), .A2(\myexu/myalu/_1016_ ), .A3(\myexu/myalu/_1018_ ), .A4(\myexu/myalu/_1019_ ), .ZN(\myexu/myalu/_1020_ ) );
OR4_X1 \myexu/myalu/_2007_ ( .A1(\myexu/myalu/_1002_ ), .A2(\myexu/myalu/_1006_ ), .A3(\myexu/myalu/_1009_ ), .A4(\myexu/myalu/_1020_ ), .ZN(\myexu/myalu/_1323_ ) );
AND3_X1 \myexu/myalu/_2008_ ( .A1(\myexu/myalu/_0687_ ), .A2(\myexu/myalu/_0773_ ), .A3(\myexu/myalu/_0905_ ), .ZN(\myexu/myalu/_1021_ ) );
AOI21_X1 \myexu/myalu/_2009_ ( .A(fanout_net_13 ), .B1(\myexu/myalu/_0854_ ), .B2(\myexu/myalu/_0856_ ), .ZN(\myexu/myalu/_1022_ ) );
AND3_X1 \myexu/myalu/_2010_ ( .A1(\myexu/myalu/_0859_ ), .A2(\myexu/myalu/_0860_ ), .A3(fanout_net_13 ), .ZN(\myexu/myalu/_1023_ ) );
NOR2_X1 \myexu/myalu/_2011_ ( .A1(\myexu/myalu/_1022_ ), .A2(\myexu/myalu/_1023_ ), .ZN(\myexu/myalu/_1024_ ) );
MUX2_X1 \myexu/myalu/_2012_ ( .A(\myexu/myalu/_1021_ ), .B(\myexu/myalu/_1024_ ), .S(\myexu/myalu/_0506_ ), .Z(\myexu/myalu/_1025_ ) );
AND2_X1 \myexu/myalu/_2013_ ( .A1(\myexu/myalu/_1025_ ), .A2(fanout_net_17 ), .ZN(\myexu/myalu/_1026_ ) );
AND2_X1 \myexu/myalu/_2014_ ( .A1(\myexu/myalu/_0845_ ), .A2(\myexu/myalu/_0846_ ), .ZN(\myexu/myalu/_1027_ ) );
MUX2_X1 \myexu/myalu/_2015_ ( .A(\myexu/myalu/_0852_ ), .B(\myexu/myalu/_1027_ ), .S(\myexu/myalu/_0703_ ), .Z(\myexu/myalu/_1028_ ) );
NAND2_X1 \myexu/myalu/_2016_ ( .A1(\myexu/myalu/_1028_ ), .A2(fanout_net_15 ), .ZN(\myexu/myalu/_1029_ ) );
NAND3_X1 \myexu/myalu/_2017_ ( .A1(\myexu/myalu/_0833_ ), .A2(\myexu/myalu/_0834_ ), .A3(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_1030_ ) );
OAI211_X2 \myexu/myalu/_2018_ ( .A(\myexu/myalu/_1030_ ), .B(\myexu/myalu/_0995_ ), .C1(\myexu/myalu/_0842_ ), .C2(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_1031_ ) );
AOI21_X1 \myexu/myalu/_2019_ ( .A(fanout_net_17 ), .B1(\myexu/myalu/_1029_ ), .B2(\myexu/myalu/_1031_ ), .ZN(\myexu/myalu/_1032_ ) );
NOR2_X1 \myexu/myalu/_2020_ ( .A1(\myexu/myalu/_1026_ ), .A2(\myexu/myalu/_1032_ ), .ZN(\myexu/myalu/_1033_ ) );
NOR2_X1 \myexu/myalu/_2021_ ( .A1(\myexu/myalu/_1033_ ), .A2(\myexu/myalu/_0734_ ), .ZN(\myexu/myalu/_1034_ ) );
AND2_X1 \myexu/myalu/_2022_ ( .A1(\myexu/myalu/_0633_ ), .A2(\myexu/myalu/_0803_ ), .ZN(\myexu/myalu/_1035_ ) );
OAI211_X2 \myexu/myalu/_2023_ ( .A(\myexu/myalu/_1035_ ), .B(\myexu/myalu/_0812_ ), .C1(fanout_net_14 ), .C2(\myexu/myalu/_0660_ ), .ZN(\myexu/myalu/_1036_ ) );
AOI21_X1 \myexu/myalu/_2024_ ( .A(\myexu/myalu/_0950_ ), .B1(\myexu/myalu/_1036_ ), .B2(\myexu/myalu/_1033_ ), .ZN(\myexu/myalu/_1037_ ) );
OAI211_X2 \myexu/myalu/_2025_ ( .A(\myexu/myalu/_0482_ ), .B(\myexu/myalu/_0491_ ), .C1(\myexu/myalu/_0967_ ), .C2(\myexu/myalu/_0969_ ), .ZN(\myexu/myalu/_1038_ ) );
AOI21_X2 \myexu/myalu/_2026_ ( .A(\myexu/myalu/_1017_ ), .B1(\myexu/myalu/_0482_ ), .B2(\myexu/myalu/_0984_ ), .ZN(\myexu/myalu/_1039_ ) );
AND2_X1 \myexu/myalu/_2027_ ( .A1(\myexu/myalu/_1038_ ), .A2(\myexu/myalu/_1039_ ), .ZN(\myexu/myalu/_1040_ ) );
INV_X1 \myexu/myalu/_2028_ ( .A(\myexu/myalu/_0487_ ), .ZN(\myexu/myalu/_1041_ ) );
OAI21_X1 \myexu/myalu/_2029_ ( .A(\myexu/myalu/_0827_ ), .B1(\myexu/myalu/_1040_ ), .B2(\myexu/myalu/_1041_ ), .ZN(\myexu/myalu/_1042_ ) );
AOI21_X1 \myexu/myalu/_2030_ ( .A(\myexu/myalu/_1042_ ), .B1(\myexu/myalu/_1041_ ), .B2(\myexu/myalu/_1040_ ), .ZN(\myexu/myalu/_1043_ ) );
OR3_X1 \myexu/myalu/_2031_ ( .A1(\myexu/myalu/_0669_ ), .A2(\myexu/myalu/_0662_ ), .A3(\myexu/myalu/_0664_ ), .ZN(\myexu/myalu/_1044_ ) );
OR3_X1 \myexu/myalu/_2032_ ( .A1(\myexu/myalu/_0666_ ), .A2(\myexu/myalu/_0670_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_1045_ ) );
AND2_X1 \myexu/myalu/_2033_ ( .A1(\myexu/myalu/_1044_ ), .A2(\myexu/myalu/_1045_ ), .ZN(\myexu/myalu/_1046_ ) );
MUX2_X1 \myexu/myalu/_2034_ ( .A(\myexu/myalu/_0879_ ), .B(\myexu/myalu/_1046_ ), .S(\myexu/myalu/_0703_ ), .Z(\myexu/myalu/_1047_ ) );
NAND3_X1 \myexu/myalu/_2035_ ( .A1(\myexu/myalu/_1047_ ), .A2(\myexu/myalu/_0980_ ), .A3(\myexu/myalu/_0885_ ), .ZN(\myexu/myalu/_1048_ ) );
NAND2_X1 \myexu/myalu/_2036_ ( .A1(\myexu/myalu/_0487_ ), .A2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_1049_ ) );
AND2_X1 \myexu/myalu/_2037_ ( .A1(\myexu/myalu/_1388_ ), .A2(\myexu/myalu/_1356_ ), .ZN(\myexu/myalu/_1050_ ) );
NAND3_X1 \myexu/myalu/_2038_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0729_ ), .A3(\myexu/myalu/_1050_ ), .ZN(\myexu/myalu/_1051_ ) );
OAI21_X1 \myexu/myalu/_2039_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1388_ ), .B2(\myexu/myalu/_1356_ ), .ZN(\myexu/myalu/_1052_ ) );
NAND4_X1 \myexu/myalu/_2040_ ( .A1(\myexu/myalu/_1048_ ), .A2(\myexu/myalu/_1049_ ), .A3(\myexu/myalu/_1051_ ), .A4(\myexu/myalu/_1052_ ), .ZN(\myexu/myalu/_1053_ ) );
OR4_X1 \myexu/myalu/_2041_ ( .A1(\myexu/myalu/_1034_ ), .A2(\myexu/myalu/_1037_ ), .A3(\myexu/myalu/_1043_ ), .A4(\myexu/myalu/_1053_ ), .ZN(\myexu/myalu/_1324_ ) );
INV_X1 \myexu/myalu/_2042_ ( .A(\myexu/myalu/_0488_ ), .ZN(\myexu/myalu/_1054_ ) );
INV_X1 \myexu/myalu/_2043_ ( .A(\myexu/myalu/_1050_ ), .ZN(\myexu/myalu/_1055_ ) );
OAI211_X2 \myexu/myalu/_2044_ ( .A(\myexu/myalu/_1054_ ), .B(\myexu/myalu/_1055_ ), .C1(\myexu/myalu/_1040_ ), .C2(\myexu/myalu/_1041_ ), .ZN(\myexu/myalu/_1056_ ) );
AOI21_X1 \myexu/myalu/_2045_ ( .A(\myexu/myalu/_1041_ ), .B1(\myexu/myalu/_1038_ ), .B2(\myexu/myalu/_1039_ ), .ZN(\myexu/myalu/_1057_ ) );
OAI21_X1 \myexu/myalu/_2046_ ( .A(\myexu/myalu/_0488_ ), .B1(\myexu/myalu/_1057_ ), .B2(\myexu/myalu/_1050_ ), .ZN(\myexu/myalu/_1058_ ) );
AND3_X1 \myexu/myalu/_2047_ ( .A1(\myexu/myalu/_1056_ ), .A2(\myexu/myalu/_0827_ ), .A3(\myexu/myalu/_1058_ ), .ZN(\myexu/myalu/_1059_ ) );
INV_X1 \myexu/myalu/_2048_ ( .A(\myexu/myalu/_0678_ ), .ZN(\myexu/myalu/_1060_ ) );
AND2_X1 \myexu/myalu/_2049_ ( .A1(\myexu/myalu/_0633_ ), .A2(\myexu/myalu/_0810_ ), .ZN(\myexu/myalu/_1061_ ) );
BUF_X4 \myexu/myalu/_2050_ ( .A(\myexu/myalu/_1061_ ), .Z(\myexu/myalu/_1062_ ) );
BUF_X2 \myexu/myalu/_2051_ ( .A(\myexu/myalu/_0811_ ), .Z(\myexu/myalu/_1063_ ) );
AND4_X1 \myexu/myalu/_2052_ ( .A1(\myexu/myalu/_1062_ ), .A2(\myexu/myalu/_0636_ ), .A3(\myexu/myalu/_1063_ ), .A4(\myexu/myalu/_0803_ ), .ZN(\myexu/myalu/_1064_ ) );
AND3_X1 \myexu/myalu/_2053_ ( .A1(\myexu/myalu/_0584_ ), .A2(\myexu/myalu/_0773_ ), .A3(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_1065_ ) );
NAND3_X1 \myexu/myalu/_2054_ ( .A1(\myexu/myalu/_0895_ ), .A2(\myexu/myalu/_0896_ ), .A3(\myexu/myalu/_0773_ ), .ZN(\myexu/myalu/_1066_ ) );
NAND3_X1 \myexu/myalu/_2055_ ( .A1(\myexu/myalu/_0902_ ), .A2(\myexu/myalu/_0903_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_1067_ ) );
NAND2_X1 \myexu/myalu/_2056_ ( .A1(\myexu/myalu/_1066_ ), .A2(\myexu/myalu/_1067_ ), .ZN(\myexu/myalu/_1068_ ) );
MUX2_X1 \myexu/myalu/_2057_ ( .A(\myexu/myalu/_1065_ ), .B(\myexu/myalu/_1068_ ), .S(\myexu/myalu/_0882_ ), .Z(\myexu/myalu/_1069_ ) );
NAND2_X1 \myexu/myalu/_2058_ ( .A1(\myexu/myalu/_1069_ ), .A2(fanout_net_17 ), .ZN(\myexu/myalu/_1070_ ) );
AOI21_X1 \myexu/myalu/_2059_ ( .A(\myexu/myalu/_0703_ ), .B1(\myexu/myalu/_0898_ ), .B2(\myexu/myalu/_0899_ ), .ZN(\myexu/myalu/_1071_ ) );
AOI21_X1 \myexu/myalu/_2060_ ( .A(fanout_net_14 ), .B1(\myexu/myalu/_0915_ ), .B2(\myexu/myalu/_0916_ ), .ZN(\myexu/myalu/_1072_ ) );
OAI21_X1 \myexu/myalu/_2061_ ( .A(fanout_net_15 ), .B1(\myexu/myalu/_1071_ ), .B2(\myexu/myalu/_1072_ ), .ZN(\myexu/myalu/_1073_ ) );
AND2_X1 \myexu/myalu/_2062_ ( .A1(\myexu/myalu/_0912_ ), .A2(\myexu/myalu/_0913_ ), .ZN(\myexu/myalu/_1074_ ) );
MUX2_X1 \myexu/myalu/_2063_ ( .A(\myexu/myalu/_0921_ ), .B(\myexu/myalu/_1074_ ), .S(fanout_net_14 ), .Z(\myexu/myalu/_1075_ ) );
OAI211_X2 \myexu/myalu/_2064_ ( .A(\myexu/myalu/_0866_ ), .B(\myexu/myalu/_1073_ ), .C1(\myexu/myalu/_1075_ ), .C2(fanout_net_15 ), .ZN(\myexu/myalu/_1076_ ) );
NAND2_X1 \myexu/myalu/_2065_ ( .A1(\myexu/myalu/_1070_ ), .A2(\myexu/myalu/_1076_ ), .ZN(\myexu/myalu/_1077_ ) );
OAI21_X1 \myexu/myalu/_2066_ ( .A(\myexu/myalu/_1060_ ), .B1(\myexu/myalu/_1064_ ), .B2(\myexu/myalu/_1077_ ), .ZN(\myexu/myalu/_1078_ ) );
OAI21_X1 \myexu/myalu/_2067_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0789_ ), .B2(\myexu/myalu/_0784_ ), .ZN(\myexu/myalu/_1079_ ) );
OAI21_X1 \myexu/myalu/_2068_ ( .A(\myexu/myalu/_0905_ ), .B1(\myexu/myalu/_0792_ ), .B2(\myexu/myalu/_0790_ ), .ZN(\myexu/myalu/_1080_ ) );
NAND2_X1 \myexu/myalu/_2069_ ( .A1(\myexu/myalu/_1079_ ), .A2(\myexu/myalu/_1080_ ), .ZN(\myexu/myalu/_1081_ ) );
NAND2_X1 \myexu/myalu/_2070_ ( .A1(\myexu/myalu/_1081_ ), .A2(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_1082_ ) );
OAI21_X1 \myexu/myalu/_2071_ ( .A(\myexu/myalu/_1082_ ), .B1(\myexu/myalu/_0940_ ), .B2(\myexu/myalu/_0843_ ), .ZN(\myexu/myalu/_1083_ ) );
NAND3_X1 \myexu/myalu/_2072_ ( .A1(\myexu/myalu/_1083_ ), .A2(\myexu/myalu/_0980_ ), .A3(\myexu/myalu/_0886_ ), .ZN(\myexu/myalu/_1084_ ) );
NAND2_X1 \myexu/myalu/_2073_ ( .A1(\myexu/myalu/_1078_ ), .A2(\myexu/myalu/_1084_ ), .ZN(\myexu/myalu/_1085_ ) );
AND3_X1 \myexu/myalu/_2074_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0478_ ), .ZN(\myexu/myalu/_1086_ ) );
NAND3_X1 \myexu/myalu/_2075_ ( .A1(\myexu/myalu/_0488_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0635_ ), .ZN(\myexu/myalu/_1087_ ) );
OAI21_X1 \myexu/myalu/_2076_ ( .A(\myexu/myalu/_1087_ ), .B1(\myexu/myalu/_0872_ ), .B2(\myexu/myalu/_0479_ ), .ZN(\myexu/myalu/_1088_ ) );
OR4_X1 \myexu/myalu/_2077_ ( .A1(\myexu/myalu/_1059_ ), .A2(\myexu/myalu/_1085_ ), .A3(\myexu/myalu/_1086_ ), .A4(\myexu/myalu/_1088_ ), .ZN(\myexu/myalu/_1325_ ) );
OR2_X1 \myexu/myalu/_2078_ ( .A1(\myexu/myalu/_0586_ ), .A2(fanout_net_15 ), .ZN(\myexu/myalu/_1089_ ) );
AND4_X1 \myexu/myalu/_2079_ ( .A1(\myexu/myalu/_0810_ ), .A2(\myexu/myalu/_0634_ ), .A3(\myexu/myalu/_1063_ ), .A4(\myexu/myalu/_1089_ ), .ZN(\myexu/myalu/_1090_ ) );
BUF_X4 \myexu/myalu/_2080_ ( .A(\myexu/myalu/_1000_ ), .Z(\myexu/myalu/_1091_ ) );
NAND3_X1 \myexu/myalu/_2081_ ( .A1(\myexu/myalu/_0693_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_1091_ ), .ZN(\myexu/myalu/_1092_ ) );
NAND3_X1 \myexu/myalu/_2082_ ( .A1(\myexu/myalu/_0647_ ), .A2(\myexu/myalu/_0654_ ), .A3(\myexu/myalu/_1000_ ), .ZN(\myexu/myalu/_1093_ ) );
OAI211_X2 \myexu/myalu/_2083_ ( .A(\myexu/myalu/_1093_ ), .B(\myexu/myalu/_0911_ ), .C1(\myexu/myalu/_0713_ ), .C2(\myexu/myalu/_1091_ ), .ZN(\myexu/myalu/_1094_ ) );
NAND2_X1 \myexu/myalu/_2084_ ( .A1(\myexu/myalu/_1092_ ), .A2(\myexu/myalu/_1094_ ), .ZN(\myexu/myalu/_1095_ ) );
OAI21_X1 \myexu/myalu/_2085_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_1090_ ), .B2(\myexu/myalu/_1095_ ), .ZN(\myexu/myalu/_1096_ ) );
NAND2_X1 \myexu/myalu/_2086_ ( .A1(\myexu/myalu/_1095_ ), .A2(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_1097_ ) );
NOR3_X2 \myexu/myalu/_2087_ ( .A1(\myexu/myalu/_1039_ ), .A2(\myexu/myalu/_1054_ ), .A3(\myexu/myalu/_1041_ ), .ZN(\myexu/myalu/_1098_ ) );
AOI211_X2 \myexu/myalu/_2088_ ( .A(\myexu/myalu/_0478_ ), .B(\myexu/myalu/_1098_ ), .C1(\myexu/myalu/_0488_ ), .C2(\myexu/myalu/_1050_ ), .ZN(\myexu/myalu/_1099_ ) );
AND4_X1 \myexu/myalu/_2089_ ( .A1(\myexu/myalu/_0488_ ), .A2(\myexu/myalu/_0487_ ), .A3(\myexu/myalu/_0482_ ), .A4(\myexu/myalu/_0491_ ), .ZN(\myexu/myalu/_1100_ ) );
OAI21_X2 \myexu/myalu/_2090_ ( .A(\myexu/myalu/_1100_ ), .B1(\myexu/myalu/_0967_ ), .B2(\myexu/myalu/_0969_ ), .ZN(\myexu/myalu/_1101_ ) );
AND2_X4 \myexu/myalu/_2091_ ( .A1(\myexu/myalu/_1099_ ), .A2(\myexu/myalu/_1101_ ), .ZN(\myexu/myalu/_1102_ ) );
AOI21_X1 \myexu/myalu/_2092_ ( .A(\myexu/myalu/_0932_ ), .B1(\myexu/myalu/_1102_ ), .B2(\myexu/myalu/_0474_ ), .ZN(\myexu/myalu/_1103_ ) );
OAI21_X1 \myexu/myalu/_2093_ ( .A(\myexu/myalu/_1103_ ), .B1(\myexu/myalu/_0474_ ), .B2(\myexu/myalu/_1102_ ), .ZN(\myexu/myalu/_1104_ ) );
NAND2_X1 \myexu/myalu/_2094_ ( .A1(\myexu/myalu/_0473_ ), .A2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_1105_ ) );
OAI21_X1 \myexu/myalu/_2095_ ( .A(\myexu/myalu/_0839_ ), .B1(\myexu/myalu/_0643_ ), .B2(\myexu/myalu/_0667_ ), .ZN(\myexu/myalu/_1106_ ) );
OAI21_X1 \myexu/myalu/_2096_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0666_ ), .B2(\myexu/myalu/_0670_ ), .ZN(\myexu/myalu/_1107_ ) );
AOI21_X1 \myexu/myalu/_2097_ ( .A(fanout_net_14 ), .B1(\myexu/myalu/_1106_ ), .B2(\myexu/myalu/_1107_ ), .ZN(\myexu/myalu/_1108_ ) );
AOI21_X1 \myexu/myalu/_2098_ ( .A(\myexu/myalu/_1108_ ), .B1(fanout_net_14 ), .B2(\myexu/myalu/_0977_ ), .ZN(\myexu/myalu/_1109_ ) );
OR2_X1 \myexu/myalu/_2099_ ( .A1(\myexu/myalu/_1109_ ), .A2(fanout_net_15 ), .ZN(\myexu/myalu/_1110_ ) );
NAND4_X1 \myexu/myalu/_2100_ ( .A1(\myexu/myalu/_0584_ ), .A2(\myexu/myalu/_1328_ ), .A3(fanout_net_15 ), .A4(\myexu/myalu/_0873_ ), .ZN(\myexu/myalu/_1111_ ) );
NAND2_X1 \myexu/myalu/_2101_ ( .A1(\myexu/myalu/_1110_ ), .A2(\myexu/myalu/_1111_ ), .ZN(\myexu/myalu/_1112_ ) );
NAND2_X1 \myexu/myalu/_2102_ ( .A1(\myexu/myalu/_1112_ ), .A2(\myexu/myalu/_0886_ ), .ZN(\myexu/myalu/_1113_ ) );
AND2_X1 \myexu/myalu/_2103_ ( .A1(\myexu/myalu/_1390_ ), .A2(\myexu/myalu/_1358_ ), .ZN(\myexu/myalu/_1114_ ) );
NAND3_X1 \myexu/myalu/_2104_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_1114_ ), .ZN(\myexu/myalu/_1115_ ) );
OAI21_X1 \myexu/myalu/_2105_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1390_ ), .B2(\myexu/myalu/_1358_ ), .ZN(\myexu/myalu/_1116_ ) );
AND4_X1 \myexu/myalu/_2106_ ( .A1(\myexu/myalu/_1105_ ), .A2(\myexu/myalu/_1113_ ), .A3(\myexu/myalu/_1115_ ), .A4(\myexu/myalu/_1116_ ), .ZN(\myexu/myalu/_1117_ ) );
NAND4_X1 \myexu/myalu/_2107_ ( .A1(\myexu/myalu/_1096_ ), .A2(\myexu/myalu/_1097_ ), .A3(\myexu/myalu/_1104_ ), .A4(\myexu/myalu/_1117_ ), .ZN(\myexu/myalu/_1326_ ) );
NAND3_X1 \myexu/myalu/_2108_ ( .A1(\myexu/myalu/_0774_ ), .A2(\myexu/myalu/_0781_ ), .A3(\myexu/myalu/_0882_ ), .ZN(\myexu/myalu/_1118_ ) );
OAI211_X2 \myexu/myalu/_2109_ ( .A(\myexu/myalu/_1118_ ), .B(\myexu/myalu/_0866_ ), .C1(\myexu/myalu/_0751_ ), .C2(\myexu/myalu/_0883_ ), .ZN(\myexu/myalu/_1119_ ) );
NAND3_X1 \myexu/myalu/_2110_ ( .A1(\myexu/myalu/_0763_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0883_ ), .ZN(\myexu/myalu/_1120_ ) );
AOI21_X1 \myexu/myalu/_2111_ ( .A(\myexu/myalu/_0734_ ), .B1(\myexu/myalu/_1119_ ), .B2(\myexu/myalu/_1120_ ), .ZN(\myexu/myalu/_1121_ ) );
NAND3_X1 \myexu/myalu/_2112_ ( .A1(\myexu/myalu/_1012_ ), .A2(\myexu/myalu/_1011_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_1122_ ) );
OR3_X1 \myexu/myalu/_2113_ ( .A1(\myexu/myalu/_0792_ ), .A2(\myexu/myalu/_0790_ ), .A3(\myexu/myalu/_0788_ ), .ZN(\myexu/myalu/_1123_ ) );
OR3_X1 \myexu/myalu/_2114_ ( .A1(\myexu/myalu/_0769_ ), .A2(\myexu/myalu/_0793_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_1124_ ) );
NAND3_X1 \myexu/myalu/_2115_ ( .A1(\myexu/myalu/_1123_ ), .A2(\myexu/myalu/_1124_ ), .A3(\myexu/myalu/_0703_ ), .ZN(\myexu/myalu/_1125_ ) );
NAND3_X1 \myexu/myalu/_2116_ ( .A1(\myexu/myalu/_1122_ ), .A2(\myexu/myalu/_1125_ ), .A3(\myexu/myalu/_0995_ ), .ZN(\myexu/myalu/_1126_ ) );
NAND2_X1 \myexu/myalu/_2117_ ( .A1(\myexu/myalu/_0800_ ), .A2(fanout_net_15 ), .ZN(\myexu/myalu/_1127_ ) );
AND3_X1 \myexu/myalu/_2118_ ( .A1(\myexu/myalu/_1126_ ), .A2(\myexu/myalu/_0885_ ), .A3(\myexu/myalu/_1127_ ), .ZN(\myexu/myalu/_1128_ ) );
NOR2_X1 \myexu/myalu/_2119_ ( .A1(\myexu/myalu/_0804_ ), .A2(\myexu/myalu/_0807_ ), .ZN(\myexu/myalu/_1129_ ) );
NOR2_X1 \myexu/myalu/_2120_ ( .A1(\myexu/myalu/_1129_ ), .A2(fanout_net_15 ), .ZN(\myexu/myalu/_1130_ ) );
INV_X1 \myexu/myalu/_2121_ ( .A(\myexu/myalu/_1130_ ), .ZN(\myexu/myalu/_1131_ ) );
AND3_X1 \myexu/myalu/_2122_ ( .A1(\myexu/myalu/_1061_ ), .A2(\myexu/myalu/_0811_ ), .A3(\myexu/myalu/_1131_ ), .ZN(\myexu/myalu/_1132_ ) );
OAI21_X1 \myexu/myalu/_2123_ ( .A(\myexu/myalu/_1132_ ), .B1(\myexu/myalu/_0660_ ), .B2(\myexu/myalu/_0803_ ), .ZN(\myexu/myalu/_1133_ ) );
NOR3_X1 \myexu/myalu/_2124_ ( .A1(\myexu/myalu/_0839_ ), .A2(\myexu/myalu/_1360_ ), .A3(fanout_net_15 ), .ZN(\myexu/myalu/_1134_ ) );
OAI211_X2 \myexu/myalu/_2125_ ( .A(\myexu/myalu/_1119_ ), .B(\myexu/myalu/_1120_ ), .C1(\myexu/myalu/_1133_ ), .C2(\myexu/myalu/_1134_ ), .ZN(\myexu/myalu/_1135_ ) );
AOI211_X2 \myexu/myalu/_2126_ ( .A(\myexu/myalu/_1121_ ), .B(\myexu/myalu/_1128_ ), .C1(\myexu/myalu/_1135_ ), .C2(\myexu/myalu/_0815_ ), .ZN(\myexu/myalu/_1136_ ) );
AOI21_X1 \myexu/myalu/_2127_ ( .A(\myexu/myalu/_0474_ ), .B1(\myexu/myalu/_1099_ ), .B2(\myexu/myalu/_1101_ ), .ZN(\myexu/myalu/_1137_ ) );
NOR2_X1 \myexu/myalu/_2128_ ( .A1(\myexu/myalu/_1137_ ), .A2(\myexu/myalu/_1114_ ), .ZN(\myexu/myalu/_1138_ ) );
AOI21_X1 \myexu/myalu/_2129_ ( .A(\myexu/myalu/_0932_ ), .B1(\myexu/myalu/_1138_ ), .B2(\myexu/myalu/_0472_ ), .ZN(\myexu/myalu/_1139_ ) );
OAI21_X1 \myexu/myalu/_2130_ ( .A(\myexu/myalu/_1139_ ), .B1(\myexu/myalu/_0472_ ), .B2(\myexu/myalu/_1138_ ), .ZN(\myexu/myalu/_1140_ ) );
NAND3_X1 \myexu/myalu/_2131_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0469_ ), .ZN(\myexu/myalu/_1141_ ) );
NOR4_X1 \myexu/myalu/_2132_ ( .A1(\myexu/myalu/_0470_ ), .A2(\myexu/myalu/_0675_ ), .A3(\myexu/myalu/_0000_ ), .A4(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_1142_ ) );
AOI21_X1 \myexu/myalu/_2133_ ( .A(\myexu/myalu/_1142_ ), .B1(\myexu/myalu/_0471_ ), .B2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_1143_ ) );
NAND4_X1 \myexu/myalu/_2134_ ( .A1(\myexu/myalu/_1136_ ), .A2(\myexu/myalu/_1140_ ), .A3(\myexu/myalu/_1141_ ), .A4(\myexu/myalu/_1143_ ), .ZN(\myexu/myalu/_1327_ ) );
INV_X1 \myexu/myalu/_2135_ ( .A(\myexu/myalu/_1132_ ), .ZN(\myexu/myalu/_1144_ ) );
AND2_X1 \myexu/myalu/_2136_ ( .A1(\myexu/myalu/_0659_ ), .A2(\myexu/myalu/_0882_ ), .ZN(\myexu/myalu/_1145_ ) );
NOR2_X1 \myexu/myalu/_2137_ ( .A1(\myexu/myalu/_1144_ ), .A2(\myexu/myalu/_1145_ ), .ZN(\myexu/myalu/_1146_ ) );
NAND3_X1 \myexu/myalu/_2138_ ( .A1(\myexu/myalu/_0853_ ), .A2(\myexu/myalu/_0857_ ), .A3(fanout_net_15 ), .ZN(\myexu/myalu/_1147_ ) );
OAI211_X2 \myexu/myalu/_2139_ ( .A(\myexu/myalu/_1147_ ), .B(\myexu/myalu/_0911_ ), .C1(\myexu/myalu/_0848_ ), .C2(fanout_net_16 ), .ZN(\myexu/myalu/_1148_ ) );
NAND3_X1 \myexu/myalu/_2140_ ( .A1(\myexu/myalu/_0863_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_1091_ ), .ZN(\myexu/myalu/_1149_ ) );
NAND2_X1 \myexu/myalu/_2141_ ( .A1(\myexu/myalu/_1148_ ), .A2(\myexu/myalu/_1149_ ), .ZN(\myexu/myalu/_1150_ ) );
OAI21_X1 \myexu/myalu/_2142_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_1146_ ), .B2(\myexu/myalu/_1150_ ), .ZN(\myexu/myalu/_1151_ ) );
INV_X1 \myexu/myalu/_2143_ ( .A(\myexu/myalu/_0464_ ), .ZN(\myexu/myalu/_1152_ ) );
AND2_X1 \myexu/myalu/_2144_ ( .A1(\myexu/myalu/_0473_ ), .A2(\myexu/myalu/_0471_ ), .ZN(\myexu/myalu/_1153_ ) );
INV_X1 \myexu/myalu/_2145_ ( .A(\myexu/myalu/_1153_ ), .ZN(\myexu/myalu/_1154_ ) );
OR2_X1 \myexu/myalu/_2146_ ( .A1(\myexu/myalu/_1102_ ), .A2(\myexu/myalu/_1154_ ), .ZN(\myexu/myalu/_1155_ ) );
AOI22_X1 \myexu/myalu/_2147_ ( .A1(\myexu/myalu/_1390_ ), .A2(\myexu/myalu/_1358_ ), .B1(\myexu/myalu/_1391_ ), .B2(\myexu/myalu/_1359_ ), .ZN(\myexu/myalu/_1156_ ) );
OR2_X4 \myexu/myalu/_2148_ ( .A1(\myexu/myalu/_1156_ ), .A2(\myexu/myalu/_0470_ ), .ZN(\myexu/myalu/_1157_ ) );
AOI21_X1 \myexu/myalu/_2149_ ( .A(\myexu/myalu/_1152_ ), .B1(\myexu/myalu/_1155_ ), .B2(\myexu/myalu/_1157_ ), .ZN(\myexu/myalu/_1158_ ) );
INV_X1 \myexu/myalu/_2150_ ( .A(\myexu/myalu/_1158_ ), .ZN(\myexu/myalu/_1159_ ) );
OAI211_X2 \myexu/myalu/_2151_ ( .A(\myexu/myalu/_1152_ ), .B(\myexu/myalu/_1157_ ), .C1(\myexu/myalu/_1102_ ), .C2(\myexu/myalu/_1154_ ), .ZN(\myexu/myalu/_1160_ ) );
NAND3_X1 \myexu/myalu/_2152_ ( .A1(\myexu/myalu/_1159_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_1160_ ), .ZN(\myexu/myalu/_1161_ ) );
NAND2_X1 \myexu/myalu/_2153_ ( .A1(\myexu/myalu/_1150_ ), .A2(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_1162_ ) );
NAND2_X1 \myexu/myalu/_2154_ ( .A1(\myexu/myalu/_0464_ ), .A2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_1163_ ) );
NAND3_X1 \myexu/myalu/_2155_ ( .A1(\myexu/myalu/_1044_ ), .A2(\myexu/myalu/_1045_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_1164_ ) );
OR3_X1 \myexu/myalu/_2156_ ( .A1(\myexu/myalu/_0643_ ), .A2(\myexu/myalu/_0667_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_1165_ ) );
OR3_X1 \myexu/myalu/_2157_ ( .A1(\myexu/myalu/_0638_ ), .A2(\myexu/myalu/_0644_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_1166_ ) );
NAND3_X1 \myexu/myalu/_2158_ ( .A1(\myexu/myalu/_1165_ ), .A2(\myexu/myalu/_1166_ ), .A3(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_1167_ ) );
NAND3_X1 \myexu/myalu/_2159_ ( .A1(\myexu/myalu/_1164_ ), .A2(\myexu/myalu/_1167_ ), .A3(\myexu/myalu/_0882_ ), .ZN(\myexu/myalu/_1168_ ) );
OAI211_X2 \myexu/myalu/_2160_ ( .A(\myexu/myalu/_1168_ ), .B(\myexu/myalu/_0910_ ), .C1(\myexu/myalu/_1000_ ), .C2(\myexu/myalu/_0881_ ), .ZN(\myexu/myalu/_1169_ ) );
OR2_X1 \myexu/myalu/_2161_ ( .A1(\myexu/myalu/_1169_ ), .A2(\myexu/myalu/_0801_ ), .ZN(\myexu/myalu/_1170_ ) );
AND2_X1 \myexu/myalu/_2162_ ( .A1(\myexu/myalu/_1361_ ), .A2(\myexu/myalu/_1329_ ), .ZN(\myexu/myalu/_1171_ ) );
NAND3_X1 \myexu/myalu/_2163_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_1171_ ), .ZN(\myexu/myalu/_1172_ ) );
OAI21_X1 \myexu/myalu/_2164_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1361_ ), .B2(\myexu/myalu/_1329_ ), .ZN(\myexu/myalu/_1173_ ) );
AND4_X1 \myexu/myalu/_2165_ ( .A1(\myexu/myalu/_1163_ ), .A2(\myexu/myalu/_1170_ ), .A3(\myexu/myalu/_1172_ ), .A4(\myexu/myalu/_1173_ ), .ZN(\myexu/myalu/_1174_ ) );
NAND4_X1 \myexu/myalu/_2166_ ( .A1(\myexu/myalu/_1151_ ), .A2(\myexu/myalu/_1161_ ), .A3(\myexu/myalu/_1162_ ), .A4(\myexu/myalu/_1174_ ), .ZN(\myexu/myalu/_1297_ ) );
OR4_X1 \myexu/myalu/_2167_ ( .A1(\myexu/myalu/_0466_ ), .A2(\myexu/myalu/_1158_ ), .A3(\myexu/myalu/_0465_ ), .A4(\myexu/myalu/_1171_ ), .ZN(\myexu/myalu/_1175_ ) );
OAI22_X1 \myexu/myalu/_2168_ ( .A1(\myexu/myalu/_1158_ ), .A2(\myexu/myalu/_1171_ ), .B1(\myexu/myalu/_0466_ ), .B2(\myexu/myalu/_0465_ ), .ZN(\myexu/myalu/_1176_ ) );
AOI21_X1 \myexu/myalu/_2169_ ( .A(\myexu/myalu/_0932_ ), .B1(\myexu/myalu/_1175_ ), .B2(\myexu/myalu/_1176_ ), .ZN(\myexu/myalu/_1177_ ) );
NAND3_X1 \myexu/myalu/_2170_ ( .A1(\myexu/myalu/_0914_ ), .A2(\myexu/myalu/_0917_ ), .A3(\myexu/myalu/_0882_ ), .ZN(\myexu/myalu/_1178_ ) );
NAND3_X1 \myexu/myalu/_2171_ ( .A1(\myexu/myalu/_0897_ ), .A2(\myexu/myalu/_0900_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_1179_ ) );
NAND3_X1 \myexu/myalu/_2172_ ( .A1(\myexu/myalu/_1178_ ), .A2(\myexu/myalu/_1179_ ), .A3(\myexu/myalu/_0865_ ), .ZN(\myexu/myalu/_1180_ ) );
AOI21_X1 \myexu/myalu/_2173_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_0904_ ), .B2(\myexu/myalu/_0906_ ), .ZN(\myexu/myalu/_1181_ ) );
NAND2_X1 \myexu/myalu/_2174_ ( .A1(\myexu/myalu/_1181_ ), .A2(fanout_net_17 ), .ZN(\myexu/myalu/_1182_ ) );
NAND2_X1 \myexu/myalu/_2175_ ( .A1(\myexu/myalu/_1180_ ), .A2(\myexu/myalu/_1182_ ), .ZN(\myexu/myalu/_1183_ ) );
OAI21_X1 \myexu/myalu/_2176_ ( .A(\myexu/myalu/_0815_ ), .B1(\myexu/myalu/_1132_ ), .B2(\myexu/myalu/_1183_ ), .ZN(\myexu/myalu/_1184_ ) );
NAND2_X1 \myexu/myalu/_2177_ ( .A1(\myexu/myalu/_1183_ ), .A2(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_1185_ ) );
OAI21_X1 \myexu/myalu/_2178_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_0940_ ), .B2(fanout_net_14 ), .ZN(\myexu/myalu/_1186_ ) );
NAND2_X1 \myexu/myalu/_2179_ ( .A1(\myexu/myalu/_1081_ ), .A2(fanout_net_14 ), .ZN(\myexu/myalu/_1187_ ) );
OR3_X1 \myexu/myalu/_2180_ ( .A1(\myexu/myalu/_0766_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0770_ ), .ZN(\myexu/myalu/_1188_ ) );
OR3_X1 \myexu/myalu/_2181_ ( .A1(\myexu/myalu/_0769_ ), .A2(\myexu/myalu/_0793_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_1189_ ) );
NAND3_X1 \myexu/myalu/_2182_ ( .A1(\myexu/myalu/_1188_ ), .A2(\myexu/myalu/_0996_ ), .A3(\myexu/myalu/_1189_ ), .ZN(\myexu/myalu/_1190_ ) );
NAND3_X1 \myexu/myalu/_2183_ ( .A1(\myexu/myalu/_1187_ ), .A2(\myexu/myalu/_1190_ ), .A3(\myexu/myalu/_1000_ ), .ZN(\myexu/myalu/_1191_ ) );
NAND3_X1 \myexu/myalu/_2184_ ( .A1(\myexu/myalu/_1186_ ), .A2(\myexu/myalu/_0885_ ), .A3(\myexu/myalu/_1191_ ), .ZN(\myexu/myalu/_1192_ ) );
NAND3_X1 \myexu/myalu/_2185_ ( .A1(\myexu/myalu/_1184_ ), .A2(\myexu/myalu/_1185_ ), .A3(\myexu/myalu/_1192_ ), .ZN(\myexu/myalu/_1193_ ) );
AND3_X1 \myexu/myalu/_2186_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0465_ ), .ZN(\myexu/myalu/_1194_ ) );
NAND3_X1 \myexu/myalu/_2187_ ( .A1(\myexu/myalu/_0467_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0635_ ), .ZN(\myexu/myalu/_1195_ ) );
OAI21_X1 \myexu/myalu/_2188_ ( .A(\myexu/myalu/_1195_ ), .B1(\myexu/myalu/_0872_ ), .B2(\myexu/myalu/_0466_ ), .ZN(\myexu/myalu/_1196_ ) );
OR4_X1 \myexu/myalu/_2189_ ( .A1(\myexu/myalu/_1177_ ), .A2(\myexu/myalu/_1193_ ), .A3(\myexu/myalu/_1194_ ), .A4(\myexu/myalu/_1196_ ), .ZN(\myexu/myalu/_1298_ ) );
OAI211_X2 \myexu/myalu/_2190_ ( .A(\myexu/myalu/_1062_ ), .B(\myexu/myalu/_1063_ ), .C1(fanout_net_16 ), .C2(\myexu/myalu/_0805_ ), .ZN(\myexu/myalu/_1197_ ) );
NOR3_X1 \myexu/myalu/_2191_ ( .A1(\myexu/myalu/_0952_ ), .A2(\myexu/myalu/_0953_ ), .A3(\myexu/myalu/_1000_ ), .ZN(\myexu/myalu/_1198_ ) );
AOI21_X1 \myexu/myalu/_2192_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_0958_ ), .B2(\myexu/myalu/_0959_ ), .ZN(\myexu/myalu/_1199_ ) );
OAI21_X1 \myexu/myalu/_2193_ ( .A(\myexu/myalu/_0867_ ), .B1(\myexu/myalu/_1198_ ), .B2(\myexu/myalu/_1199_ ), .ZN(\myexu/myalu/_1200_ ) );
NAND4_X1 \myexu/myalu/_2194_ ( .A1(\myexu/myalu/_0692_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0980_ ), .A4(\myexu/myalu/_0873_ ), .ZN(\myexu/myalu/_1201_ ) );
NAND3_X1 \myexu/myalu/_2195_ ( .A1(\myexu/myalu/_1197_ ), .A2(\myexu/myalu/_1200_ ), .A3(\myexu/myalu/_1201_ ), .ZN(\myexu/myalu/_1202_ ) );
AOI21_X1 \myexu/myalu/_2196_ ( .A(\myexu/myalu/_0734_ ), .B1(\myexu/myalu/_1200_ ), .B2(\myexu/myalu/_1201_ ), .ZN(\myexu/myalu/_1203_ ) );
OAI21_X1 \myexu/myalu/_2197_ ( .A(\myexu/myalu/_1202_ ), .B1(\myexu/myalu/_0830_ ), .B2(\myexu/myalu/_1203_ ), .ZN(\myexu/myalu/_1204_ ) );
INV_X1 \myexu/myalu/_2198_ ( .A(\myexu/myalu/_1102_ ), .ZN(\myexu/myalu/_1205_ ) );
AND2_X1 \myexu/myalu/_2199_ ( .A1(\myexu/myalu/_0464_ ), .A2(\myexu/myalu/_0467_ ), .ZN(\myexu/myalu/_1206_ ) );
AND2_X1 \myexu/myalu/_2200_ ( .A1(\myexu/myalu/_1153_ ), .A2(\myexu/myalu/_1206_ ), .ZN(\myexu/myalu/_1207_ ) );
NAND2_X1 \myexu/myalu/_2201_ ( .A1(\myexu/myalu/_1205_ ), .A2(\myexu/myalu/_1207_ ), .ZN(\myexu/myalu/_1208_ ) );
OR4_X2 \myexu/myalu/_2202_ ( .A1(\myexu/myalu/_0466_ ), .A2(\myexu/myalu/_1152_ ), .A3(\myexu/myalu/_1157_ ), .A4(\myexu/myalu/_0465_ ), .ZN(\myexu/myalu/_1209_ ) );
AOI21_X1 \myexu/myalu/_2203_ ( .A(\myexu/myalu/_0465_ ), .B1(\myexu/myalu/_0467_ ), .B2(\myexu/myalu/_1171_ ), .ZN(\myexu/myalu/_1210_ ) );
AND2_X1 \myexu/myalu/_2204_ ( .A1(\myexu/myalu/_1209_ ), .A2(\myexu/myalu/_1210_ ), .ZN(\myexu/myalu/_1211_ ) );
AND3_X1 \myexu/myalu/_2205_ ( .A1(\myexu/myalu/_1208_ ), .A2(\myexu/myalu/_0462_ ), .A3(\myexu/myalu/_1211_ ), .ZN(\myexu/myalu/_1212_ ) );
AOI21_X1 \myexu/myalu/_2206_ ( .A(\myexu/myalu/_0462_ ), .B1(\myexu/myalu/_1208_ ), .B2(\myexu/myalu/_1211_ ), .ZN(\myexu/myalu/_1213_ ) );
OR3_X1 \myexu/myalu/_2207_ ( .A1(\myexu/myalu/_1212_ ), .A2(\myexu/myalu/_1213_ ), .A3(\myexu/myalu/_0932_ ), .ZN(\myexu/myalu/_1214_ ) );
OAI21_X1 \myexu/myalu/_2208_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1363_ ), .B2(\myexu/myalu/_1331_ ), .ZN(\myexu/myalu/_1215_ ) );
NAND2_X1 \myexu/myalu/_2209_ ( .A1(\myexu/myalu/_0461_ ), .A2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_1216_ ) );
AND2_X1 \myexu/myalu/_2210_ ( .A1(\myexu/myalu/_1363_ ), .A2(\myexu/myalu/_1331_ ), .ZN(\myexu/myalu/_1217_ ) );
NAND3_X1 \myexu/myalu/_2211_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_1217_ ), .ZN(\myexu/myalu/_1218_ ) );
AND3_X1 \myexu/myalu/_2212_ ( .A1(\myexu/myalu/_1215_ ), .A2(\myexu/myalu/_1216_ ), .A3(\myexu/myalu/_1218_ ), .ZN(\myexu/myalu/_1219_ ) );
NAND2_X1 \myexu/myalu/_2213_ ( .A1(\myexu/myalu/_0979_ ), .A2(fanout_net_16 ), .ZN(\myexu/myalu/_1220_ ) );
OR3_X1 \myexu/myalu/_2214_ ( .A1(\myexu/myalu/_0638_ ), .A2(\myexu/myalu/_0644_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_1221_ ) );
OR3_X1 \myexu/myalu/_2215_ ( .A1(\myexu/myalu/_0651_ ), .A2(\myexu/myalu/_0639_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_1222_ ) );
AOI21_X1 \myexu/myalu/_2216_ ( .A(fanout_net_14 ), .B1(\myexu/myalu/_1221_ ), .B2(\myexu/myalu/_1222_ ), .ZN(\myexu/myalu/_1223_ ) );
AND3_X1 \myexu/myalu/_2217_ ( .A1(\myexu/myalu/_1106_ ), .A2(\myexu/myalu/_1107_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_1224_ ) );
OR3_X1 \myexu/myalu/_2218_ ( .A1(\myexu/myalu/_1223_ ), .A2(\myexu/myalu/_1224_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_1225_ ) );
NAND2_X1 \myexu/myalu/_2219_ ( .A1(\myexu/myalu/_1220_ ), .A2(\myexu/myalu/_1225_ ), .ZN(\myexu/myalu/_1226_ ) );
NAND2_X1 \myexu/myalu/_2220_ ( .A1(\myexu/myalu/_1226_ ), .A2(\myexu/myalu/_0886_ ), .ZN(\myexu/myalu/_1227_ ) );
NAND4_X1 \myexu/myalu/_2221_ ( .A1(\myexu/myalu/_1204_ ), .A2(\myexu/myalu/_1214_ ), .A3(\myexu/myalu/_1219_ ), .A4(\myexu/myalu/_1227_ ), .ZN(\myexu/myalu/_1299_ ) );
OR3_X1 \myexu/myalu/_2222_ ( .A1(\myexu/myalu/_1213_ ), .A2(\myexu/myalu/_0460_ ), .A3(\myexu/myalu/_1217_ ), .ZN(\myexu/myalu/_1228_ ) );
OAI21_X1 \myexu/myalu/_2223_ ( .A(\myexu/myalu/_0460_ ), .B1(\myexu/myalu/_1213_ ), .B2(\myexu/myalu/_1217_ ), .ZN(\myexu/myalu/_1229_ ) );
AOI21_X1 \myexu/myalu/_2224_ ( .A(\myexu/myalu/_0932_ ), .B1(\myexu/myalu/_1228_ ), .B2(\myexu/myalu/_1229_ ), .ZN(\myexu/myalu/_1230_ ) );
OAI211_X2 \myexu/myalu/_2225_ ( .A(\myexu/myalu/_0634_ ), .B(\myexu/myalu/_0812_ ), .C1(\myexu/myalu/_0803_ ), .C2(\myexu/myalu/_1003_ ), .ZN(\myexu/myalu/_1231_ ) );
INV_X1 \myexu/myalu/_2226_ ( .A(\myexu/myalu/_1231_ ), .ZN(\myexu/myalu/_1232_ ) );
AND3_X1 \myexu/myalu/_2227_ ( .A1(\myexu/myalu/_0989_ ), .A2(\myexu/myalu/_0990_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_1233_ ) );
AOI211_X4 \myexu/myalu/_2228_ ( .A(fanout_net_17 ), .B(\myexu/myalu/_1233_ ), .C1(\myexu/myalu/_0506_ ), .C2(\myexu/myalu/_0999_ ), .ZN(\myexu/myalu/_1234_ ) );
AND4_X1 \myexu/myalu/_2229_ ( .A1(fanout_net_17 ), .A2(\myexu/myalu/_0755_ ), .A3(\myexu/myalu/_0506_ ), .A4(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_1235_ ) );
OR2_X1 \myexu/myalu/_2230_ ( .A1(\myexu/myalu/_1234_ ), .A2(\myexu/myalu/_1235_ ), .ZN(\myexu/myalu/_1236_ ) );
OAI21_X1 \myexu/myalu/_2231_ ( .A(\myexu/myalu/_0815_ ), .B1(\myexu/myalu/_1232_ ), .B2(\myexu/myalu/_1236_ ), .ZN(\myexu/myalu/_1237_ ) );
OAI21_X1 \myexu/myalu/_2232_ ( .A(\myexu/myalu/_0929_ ), .B1(\myexu/myalu/_1234_ ), .B2(\myexu/myalu/_1235_ ), .ZN(\myexu/myalu/_1238_ ) );
AND2_X1 \myexu/myalu/_2233_ ( .A1(\myexu/myalu/_1014_ ), .A2(fanout_net_16 ), .ZN(\myexu/myalu/_1239_ ) );
OAI21_X1 \myexu/myalu/_2234_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0766_ ), .B2(\myexu/myalu/_0770_ ), .ZN(\myexu/myalu/_1240_ ) );
OAI21_X1 \myexu/myalu/_2235_ ( .A(\myexu/myalu/_0905_ ), .B1(\myexu/myalu/_0778_ ), .B2(\myexu/myalu/_0767_ ), .ZN(\myexu/myalu/_1241_ ) );
NAND2_X1 \myexu/myalu/_2236_ ( .A1(\myexu/myalu/_1240_ ), .A2(\myexu/myalu/_1241_ ), .ZN(\myexu/myalu/_1242_ ) );
NAND2_X1 \myexu/myalu/_2237_ ( .A1(\myexu/myalu/_1242_ ), .A2(\myexu/myalu/_0843_ ), .ZN(\myexu/myalu/_1243_ ) );
NAND3_X1 \myexu/myalu/_2238_ ( .A1(\myexu/myalu/_1123_ ), .A2(\myexu/myalu/_1124_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_1244_ ) );
AOI21_X1 \myexu/myalu/_2239_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_1243_ ), .B2(\myexu/myalu/_1244_ ), .ZN(\myexu/myalu/_1245_ ) );
OAI21_X1 \myexu/myalu/_2240_ ( .A(\myexu/myalu/_0885_ ), .B1(\myexu/myalu/_1239_ ), .B2(\myexu/myalu/_1245_ ), .ZN(\myexu/myalu/_1246_ ) );
NAND3_X1 \myexu/myalu/_2241_ ( .A1(\myexu/myalu/_1237_ ), .A2(\myexu/myalu/_1238_ ), .A3(\myexu/myalu/_1246_ ), .ZN(\myexu/myalu/_1247_ ) );
AND3_X1 \myexu/myalu/_2242_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0457_ ), .ZN(\myexu/myalu/_1248_ ) );
NAND3_X1 \myexu/myalu/_2243_ ( .A1(\myexu/myalu/_0459_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0635_ ), .ZN(\myexu/myalu/_1249_ ) );
OAI21_X1 \myexu/myalu/_2244_ ( .A(\myexu/myalu/_1249_ ), .B1(\myexu/myalu/_0872_ ), .B2(\myexu/myalu/_0458_ ), .ZN(\myexu/myalu/_1250_ ) );
OR4_X1 \myexu/myalu/_2245_ ( .A1(\myexu/myalu/_1230_ ), .A2(\myexu/myalu/_1247_ ), .A3(\myexu/myalu/_1248_ ), .A4(\myexu/myalu/_1250_ ), .ZN(\myexu/myalu/_1300_ ) );
AND2_X1 \myexu/myalu/_2246_ ( .A1(\myexu/myalu/_1208_ ), .A2(\myexu/myalu/_1211_ ), .ZN(\myexu/myalu/_1251_ ) );
AND2_X1 \myexu/myalu/_2247_ ( .A1(\myexu/myalu/_0461_ ), .A2(\myexu/myalu/_0459_ ), .ZN(\myexu/myalu/_1252_ ) );
INV_X1 \myexu/myalu/_2248_ ( .A(\myexu/myalu/_1252_ ), .ZN(\myexu/myalu/_1253_ ) );
OR2_X1 \myexu/myalu/_2249_ ( .A1(\myexu/myalu/_1251_ ), .A2(\myexu/myalu/_1253_ ), .ZN(\myexu/myalu/_1254_ ) );
INV_X1 \myexu/myalu/_2250_ ( .A(\myexu/myalu/_0438_ ), .ZN(\myexu/myalu/_1255_ ) );
AOI21_X1 \myexu/myalu/_2251_ ( .A(\myexu/myalu/_0457_ ), .B1(\myexu/myalu/_0459_ ), .B2(\myexu/myalu/_1217_ ), .ZN(\myexu/myalu/_1256_ ) );
AND3_X1 \myexu/myalu/_2252_ ( .A1(\myexu/myalu/_1254_ ), .A2(\myexu/myalu/_1255_ ), .A3(\myexu/myalu/_1256_ ), .ZN(\myexu/myalu/_1257_ ) );
AOI21_X1 \myexu/myalu/_2253_ ( .A(\myexu/myalu/_1255_ ), .B1(\myexu/myalu/_1254_ ), .B2(\myexu/myalu/_1256_ ), .ZN(\myexu/myalu/_1258_ ) );
NOR3_X1 \myexu/myalu/_2254_ ( .A1(\myexu/myalu/_1257_ ), .A2(\myexu/myalu/_1258_ ), .A3(\myexu/myalu/_0932_ ), .ZN(\myexu/myalu/_1259_ ) );
INV_X4 \myexu/myalu/_2255_ ( .A(\myexu/myalu/_1062_ ), .ZN(\myexu/myalu/_1260_ ) );
INV_X1 \myexu/myalu/_2256_ ( .A(\myexu/myalu/_0811_ ), .ZN(\myexu/myalu/_1261_ ) );
AND3_X1 \myexu/myalu/_2257_ ( .A1(\myexu/myalu/_0659_ ), .A2(\myexu/myalu/_0882_ ), .A3(\myexu/myalu/_0843_ ), .ZN(\myexu/myalu/_1262_ ) );
NOR3_X1 \myexu/myalu/_2258_ ( .A1(\myexu/myalu/_1260_ ), .A2(\myexu/myalu/_1261_ ), .A3(\myexu/myalu/_1262_ ), .ZN(\myexu/myalu/_1263_ ) );
OAI21_X1 \myexu/myalu/_2259_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_1022_ ), .B2(\myexu/myalu/_1023_ ), .ZN(\myexu/myalu/_1264_ ) );
OAI211_X2 \myexu/myalu/_2260_ ( .A(\myexu/myalu/_0865_ ), .B(\myexu/myalu/_1264_ ), .C1(\myexu/myalu/_1028_ ), .C2(fanout_net_16 ), .ZN(\myexu/myalu/_1265_ ) );
NAND4_X1 \myexu/myalu/_2261_ ( .A1(\myexu/myalu/_0862_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0995_ ), .A4(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_1266_ ) );
NAND2_X1 \myexu/myalu/_2262_ ( .A1(\myexu/myalu/_1265_ ), .A2(\myexu/myalu/_1266_ ), .ZN(\myexu/myalu/_1267_ ) );
OAI21_X1 \myexu/myalu/_2263_ ( .A(\myexu/myalu/_0636_ ), .B1(\myexu/myalu/_1263_ ), .B2(\myexu/myalu/_1267_ ), .ZN(\myexu/myalu/_1268_ ) );
NAND2_X1 \myexu/myalu/_2264_ ( .A1(\myexu/myalu/_1267_ ), .A2(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_1269_ ) );
AND2_X1 \myexu/myalu/_2265_ ( .A1(\myexu/myalu/_1047_ ), .A2(fanout_net_16 ), .ZN(\myexu/myalu/_1270_ ) );
OR3_X1 \myexu/myalu/_2266_ ( .A1(\myexu/myalu/_0651_ ), .A2(\myexu/myalu/_0639_ ), .A3(\myexu/myalu/_0905_ ), .ZN(\myexu/myalu/_1271_ ) );
OR3_X1 \myexu/myalu/_2267_ ( .A1(\myexu/myalu/_0648_ ), .A2(\myexu/myalu/_0652_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_1272_ ) );
NAND3_X1 \myexu/myalu/_2268_ ( .A1(\myexu/myalu/_1271_ ), .A2(\myexu/myalu/_1272_ ), .A3(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_1273_ ) );
NAND3_X1 \myexu/myalu/_2269_ ( .A1(\myexu/myalu/_1165_ ), .A2(\myexu/myalu/_1166_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_1274_ ) );
AOI21_X1 \myexu/myalu/_2270_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_1273_ ), .B2(\myexu/myalu/_1274_ ), .ZN(\myexu/myalu/_1275_ ) );
OAI21_X1 \myexu/myalu/_2271_ ( .A(\myexu/myalu/_0885_ ), .B1(\myexu/myalu/_1270_ ), .B2(\myexu/myalu/_1275_ ), .ZN(\myexu/myalu/_1276_ ) );
NAND3_X1 \myexu/myalu/_2272_ ( .A1(\myexu/myalu/_1268_ ), .A2(\myexu/myalu/_1269_ ), .A3(\myexu/myalu/_1276_ ), .ZN(\myexu/myalu/_1277_ ) );
AND2_X1 \myexu/myalu/_2273_ ( .A1(\myexu/myalu/_1365_ ), .A2(\myexu/myalu/_1333_ ), .ZN(\myexu/myalu/_1278_ ) );
AND3_X1 \myexu/myalu/_2274_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_1278_ ), .ZN(\myexu/myalu/_1279_ ) );
OAI21_X1 \myexu/myalu/_2275_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1365_ ), .B2(\myexu/myalu/_1333_ ), .ZN(\myexu/myalu/_1280_ ) );
OAI21_X1 \myexu/myalu/_2276_ ( .A(\myexu/myalu/_1280_ ), .B1(\myexu/myalu/_1255_ ), .B2(\myexu/myalu/_0722_ ), .ZN(\myexu/myalu/_1281_ ) );
OR4_X1 \myexu/myalu/_2277_ ( .A1(\myexu/myalu/_1259_ ), .A2(\myexu/myalu/_1277_ ), .A3(\myexu/myalu/_1279_ ), .A4(\myexu/myalu/_1281_ ), .ZN(\myexu/myalu/_1301_ ) );
NAND4_X1 \myexu/myalu/_2278_ ( .A1(\myexu/myalu/_0634_ ), .A2(\myexu/myalu/_0810_ ), .A3(\myexu/myalu/_0815_ ), .A4(\myexu/myalu/_1063_ ), .ZN(\myexu/myalu/_1282_ ) );
NAND4_X1 \myexu/myalu/_2279_ ( .A1(\myexu/myalu/_0586_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_1091_ ), .A4(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_1283_ ) );
OAI21_X1 \myexu/myalu/_2280_ ( .A(\myexu/myalu/_0980_ ), .B1(\myexu/myalu/_1071_ ), .B2(\myexu/myalu/_1072_ ), .ZN(\myexu/myalu/_1284_ ) );
OAI211_X2 \myexu/myalu/_2281_ ( .A(\myexu/myalu/_1284_ ), .B(\myexu/myalu/_0911_ ), .C1(\myexu/myalu/_1091_ ), .C2(\myexu/myalu/_1068_ ), .ZN(\myexu/myalu/_1285_ ) );
NAND3_X1 \myexu/myalu/_2282_ ( .A1(\myexu/myalu/_1282_ ), .A2(\myexu/myalu/_1283_ ), .A3(\myexu/myalu/_1285_ ), .ZN(\myexu/myalu/_1286_ ) );
AND2_X1 \myexu/myalu/_2283_ ( .A1(\myexu/myalu/_1083_ ), .A2(fanout_net_16 ), .ZN(\myexu/myalu/_1287_ ) );
OR3_X1 \myexu/myalu/_2284_ ( .A1(\myexu/myalu/_0775_ ), .A2(fanout_net_12 ), .A3(\myexu/myalu/_0779_ ), .ZN(\myexu/myalu/_1288_ ) );
OR3_X1 \myexu/myalu/_2285_ ( .A1(\myexu/myalu/_0778_ ), .A2(\myexu/myalu/_0767_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_1289_ ) );
NAND3_X1 \myexu/myalu/_2286_ ( .A1(\myexu/myalu/_1288_ ), .A2(\myexu/myalu/_0843_ ), .A3(\myexu/myalu/_1289_ ), .ZN(\myexu/myalu/_1290_ ) );
NAND3_X1 \myexu/myalu/_2287_ ( .A1(\myexu/myalu/_1188_ ), .A2(fanout_net_14 ), .A3(\myexu/myalu/_1189_ ), .ZN(\myexu/myalu/_1291_ ) );
AOI21_X1 \myexu/myalu/_2288_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_1290_ ), .B2(\myexu/myalu/_1291_ ), .ZN(\myexu/myalu/_1292_ ) );
OR2_X1 \myexu/myalu/_2289_ ( .A1(\myexu/myalu/_1287_ ), .A2(\myexu/myalu/_1292_ ), .ZN(\myexu/myalu/_1293_ ) );
AOI22_X1 \myexu/myalu/_2290_ ( .A1(\myexu/myalu/_1286_ ), .A2(\myexu/myalu/_1060_ ), .B1(\myexu/myalu/_0886_ ), .B2(\myexu/myalu/_1293_ ), .ZN(\myexu/myalu/_1294_ ) );
OR3_X1 \myexu/myalu/_2291_ ( .A1(\myexu/myalu/_1258_ ), .A2(\myexu/myalu/_0455_ ), .A3(\myexu/myalu/_1278_ ), .ZN(\myexu/myalu/_1295_ ) );
OAI21_X1 \myexu/myalu/_2292_ ( .A(\myexu/myalu/_0455_ ), .B1(\myexu/myalu/_1258_ ), .B2(\myexu/myalu/_1278_ ), .ZN(\myexu/myalu/_0004_ ) );
NAND3_X1 \myexu/myalu/_2293_ ( .A1(\myexu/myalu/_1295_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_0004_ ), .ZN(\myexu/myalu/_0005_ ) );
NOR4_X1 \myexu/myalu/_2294_ ( .A1(\myexu/myalu/_0454_ ), .A2(\myexu/myalu/_0675_ ), .A3(\myexu/myalu/_0000_ ), .A4(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0006_ ) );
AOI21_X1 \myexu/myalu/_2295_ ( .A(\myexu/myalu/_0006_ ), .B1(\myexu/myalu/_0455_ ), .B2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_0007_ ) );
NAND3_X1 \myexu/myalu/_2296_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0449_ ), .ZN(\myexu/myalu/_0008_ ) );
NAND4_X1 \myexu/myalu/_2297_ ( .A1(\myexu/myalu/_1294_ ), .A2(\myexu/myalu/_0005_ ), .A3(\myexu/myalu/_0007_ ), .A4(\myexu/myalu/_0008_ ), .ZN(\myexu/myalu/_1302_ ) );
INV_X1 \myexu/myalu/_2298_ ( .A(\myexu/myalu/_0417_ ), .ZN(\myexu/myalu/_0009_ ) );
NAND2_X1 \myexu/myalu/_2299_ ( .A1(\myexu/myalu/_0438_ ), .A2(\myexu/myalu/_0455_ ), .ZN(\myexu/myalu/_0010_ ) );
NOR3_X1 \myexu/myalu/_2300_ ( .A1(\myexu/myalu/_0010_ ), .A2(\myexu/myalu/_0462_ ), .A3(\myexu/myalu/_0460_ ), .ZN(\myexu/myalu/_0011_ ) );
NAND3_X2 \myexu/myalu/_2301_ ( .A1(\myexu/myalu/_1205_ ), .A2(\myexu/myalu/_1207_ ), .A3(\myexu/myalu/_0011_ ), .ZN(\myexu/myalu/_0012_ ) );
AOI211_X4 \myexu/myalu/_2302_ ( .A(\myexu/myalu/_0010_ ), .B(\myexu/myalu/_1253_ ), .C1(\myexu/myalu/_1209_ ), .C2(\myexu/myalu/_1210_ ), .ZN(\myexu/myalu/_0014_ ) );
NOR2_X1 \myexu/myalu/_2303_ ( .A1(\myexu/myalu/_1256_ ), .A2(\myexu/myalu/_0010_ ), .ZN(\myexu/myalu/_0015_ ) );
AND2_X1 \myexu/myalu/_2304_ ( .A1(\myexu/myalu/_0455_ ), .A2(\myexu/myalu/_1278_ ), .ZN(\myexu/myalu/_0016_ ) );
NOR4_X1 \myexu/myalu/_2305_ ( .A1(\myexu/myalu/_0014_ ), .A2(\myexu/myalu/_0449_ ), .A3(\myexu/myalu/_0015_ ), .A4(\myexu/myalu/_0016_ ), .ZN(\myexu/myalu/_0017_ ) );
AOI21_X1 \myexu/myalu/_2306_ ( .A(\myexu/myalu/_0009_ ), .B1(\myexu/myalu/_0012_ ), .B2(\myexu/myalu/_0017_ ), .ZN(\myexu/myalu/_0018_ ) );
INV_X1 \myexu/myalu/_2307_ ( .A(\myexu/myalu/_0018_ ), .ZN(\myexu/myalu/_0019_ ) );
NAND3_X1 \myexu/myalu/_2308_ ( .A1(\myexu/myalu/_0012_ ), .A2(\myexu/myalu/_0009_ ), .A3(\myexu/myalu/_0017_ ), .ZN(\myexu/myalu/_0020_ ) );
AND3_X1 \myexu/myalu/_2309_ ( .A1(\myexu/myalu/_0019_ ), .A2(\myexu/myalu/_0827_ ), .A3(\myexu/myalu/_0020_ ), .ZN(\myexu/myalu/_0021_ ) );
OAI211_X2 \myexu/myalu/_2310_ ( .A(\myexu/myalu/_0634_ ), .B(\myexu/myalu/_0810_ ), .C1(fanout_net_17 ), .C2(\myexu/myalu/_0587_ ), .ZN(\myexu/myalu/_0022_ ) );
OAI21_X1 \myexu/myalu/_2311_ ( .A(\myexu/myalu/_0022_ ), .B1(fanout_net_17 ), .B2(\myexu/myalu/_0714_ ), .ZN(\myexu/myalu/_0023_ ) );
AND2_X1 \myexu/myalu/_2312_ ( .A1(\myexu/myalu/_0023_ ), .A2(\myexu/myalu/_0815_ ), .ZN(\myexu/myalu/_0025_ ) );
NOR2_X1 \myexu/myalu/_2313_ ( .A1(\myexu/myalu/_1109_ ), .A2(\myexu/myalu/_1000_ ), .ZN(\myexu/myalu/_0026_ ) );
OR3_X1 \myexu/myalu/_2314_ ( .A1(\myexu/myalu/_0648_ ), .A2(\myexu/myalu/_0652_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_0027_ ) );
OR3_X1 \myexu/myalu/_2315_ ( .A1(\myexu/myalu/_0696_ ), .A2(\myexu/myalu/_0649_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0028_ ) );
NAND3_X1 \myexu/myalu/_2316_ ( .A1(\myexu/myalu/_0027_ ), .A2(\myexu/myalu/_0028_ ), .A3(\myexu/myalu/_0880_ ), .ZN(\myexu/myalu/_0029_ ) );
NAND3_X1 \myexu/myalu/_2317_ ( .A1(\myexu/myalu/_1221_ ), .A2(\myexu/myalu/_1222_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_0030_ ) );
AOI21_X1 \myexu/myalu/_2318_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_0029_ ), .B2(\myexu/myalu/_0030_ ), .ZN(\myexu/myalu/_0031_ ) );
OAI21_X1 \myexu/myalu/_2319_ ( .A(\myexu/myalu/_0867_ ), .B1(\myexu/myalu/_0026_ ), .B2(\myexu/myalu/_0031_ ), .ZN(\myexu/myalu/_0032_ ) );
NAND4_X1 \myexu/myalu/_2320_ ( .A1(\myexu/myalu/_0586_ ), .A2(\myexu/myalu/_1328_ ), .A3(fanout_net_17 ), .A4(\myexu/myalu/_0980_ ), .ZN(\myexu/myalu/_0033_ ) );
AOI21_X1 \myexu/myalu/_2321_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0032_ ), .B2(\myexu/myalu/_0033_ ), .ZN(\myexu/myalu/_0034_ ) );
OR3_X1 \myexu/myalu/_2322_ ( .A1(\myexu/myalu/_0714_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0734_ ), .ZN(\myexu/myalu/_0036_ ) );
OAI211_X2 \myexu/myalu/_2323_ ( .A(\myexu/myalu/_0676_ ), .B(\myexu/myalu/_0729_ ), .C1(\myexu/myalu/_1367_ ), .C2(\myexu/myalu/_1335_ ), .ZN(\myexu/myalu/_0037_ ) );
NAND2_X1 \myexu/myalu/_2324_ ( .A1(\myexu/myalu/_0417_ ), .A2(\myexu/myalu/_0721_ ), .ZN(\myexu/myalu/_0038_ ) );
AND2_X1 \myexu/myalu/_2325_ ( .A1(\myexu/myalu/_1367_ ), .A2(\myexu/myalu/_1335_ ), .ZN(\myexu/myalu/_0039_ ) );
NAND3_X1 \myexu/myalu/_2326_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0729_ ), .A3(\myexu/myalu/_0039_ ), .ZN(\myexu/myalu/_0040_ ) );
NAND4_X1 \myexu/myalu/_2327_ ( .A1(\myexu/myalu/_0036_ ), .A2(\myexu/myalu/_0037_ ), .A3(\myexu/myalu/_0038_ ), .A4(\myexu/myalu/_0040_ ), .ZN(\myexu/myalu/_0041_ ) );
OR4_X1 \myexu/myalu/_2328_ ( .A1(\myexu/myalu/_0021_ ), .A2(\myexu/myalu/_0025_ ), .A3(\myexu/myalu/_0034_ ), .A4(\myexu/myalu/_0041_ ), .ZN(\myexu/myalu/_1303_ ) );
NOR2_X1 \myexu/myalu/_2329_ ( .A1(\myexu/myalu/_0018_ ), .A2(\myexu/myalu/_0039_ ), .ZN(\myexu/myalu/_0042_ ) );
XNOR2_X1 \myexu/myalu/_2330_ ( .A(\myexu/myalu/_0042_ ), .B(\myexu/myalu/_0407_ ), .ZN(\myexu/myalu/_0043_ ) );
AND3_X1 \myexu/myalu/_2331_ ( .A1(\myexu/myalu/_0043_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0559_ ), .ZN(\myexu/myalu/_0044_ ) );
NOR2_X1 \myexu/myalu/_2332_ ( .A1(\myexu/myalu/_0811_ ), .A2(\myexu/myalu/_1387_ ), .ZN(\myexu/myalu/_0046_ ) );
NAND3_X1 \myexu/myalu/_2333_ ( .A1(\myexu/myalu/_0808_ ), .A2(\myexu/myalu/_0809_ ), .A3(\myexu/myalu/_0046_ ), .ZN(\myexu/myalu/_0047_ ) );
AOI22_X1 \myexu/myalu/_2334_ ( .A1(\myexu/myalu/_1062_ ), .A2(\myexu/myalu/_1063_ ), .B1(\myexu/myalu/_0865_ ), .B2(\myexu/myalu/_0764_ ), .ZN(\myexu/myalu/_0048_ ) );
AOI21_X1 \myexu/myalu/_2335_ ( .A(\myexu/myalu/_0950_ ), .B1(\myexu/myalu/_0047_ ), .B2(\myexu/myalu/_0048_ ), .ZN(\myexu/myalu/_0049_ ) );
AND3_X1 \myexu/myalu/_2336_ ( .A1(\myexu/myalu/_0764_ ), .A2(\myexu/myalu/_0865_ ), .A3(\myexu/myalu/_0677_ ), .ZN(\myexu/myalu/_0050_ ) );
NAND2_X1 \myexu/myalu/_2337_ ( .A1(\myexu/myalu/_1242_ ), .A2(fanout_net_14 ), .ZN(\myexu/myalu/_0051_ ) );
OR3_X1 \myexu/myalu/_2338_ ( .A1(\myexu/myalu/_0775_ ), .A2(\myexu/myalu/_0788_ ), .A3(\myexu/myalu/_0779_ ), .ZN(\myexu/myalu/_0052_ ) );
OR3_X1 \myexu/myalu/_2339_ ( .A1(\myexu/myalu/_0738_ ), .A2(\myexu/myalu/_0776_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0053_ ) );
NAND3_X1 \myexu/myalu/_2340_ ( .A1(\myexu/myalu/_0052_ ), .A2(\myexu/myalu/_0880_ ), .A3(\myexu/myalu/_0053_ ), .ZN(\myexu/myalu/_0054_ ) );
NAND3_X1 \myexu/myalu/_2341_ ( .A1(\myexu/myalu/_0051_ ), .A2(\myexu/myalu/_0054_ ), .A3(\myexu/myalu/_0882_ ), .ZN(\myexu/myalu/_0055_ ) );
NAND3_X1 \myexu/myalu/_2342_ ( .A1(\myexu/myalu/_1122_ ), .A2(\myexu/myalu/_1125_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_0057_ ) );
NAND3_X1 \myexu/myalu/_2343_ ( .A1(\myexu/myalu/_0055_ ), .A2(\myexu/myalu/_0057_ ), .A3(\myexu/myalu/_0865_ ), .ZN(\myexu/myalu/_0058_ ) );
NAND4_X1 \myexu/myalu/_2344_ ( .A1(\myexu/myalu/_1010_ ), .A2(fanout_net_17 ), .A3(\myexu/myalu/_0882_ ), .A4(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_0059_ ) );
AOI21_X1 \myexu/myalu/_2345_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0058_ ), .B2(\myexu/myalu/_0059_ ), .ZN(\myexu/myalu/_0060_ ) );
OR3_X1 \myexu/myalu/_2346_ ( .A1(\myexu/myalu/_0049_ ), .A2(\myexu/myalu/_0050_ ), .A3(\myexu/myalu/_0060_ ), .ZN(\myexu/myalu/_0061_ ) );
NAND3_X1 \myexu/myalu/_2347_ ( .A1(\myexu/myalu/_0407_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0635_ ), .ZN(\myexu/myalu/_0062_ ) );
OAI21_X1 \myexu/myalu/_2348_ ( .A(\myexu/myalu/_0062_ ), .B1(\myexu/myalu/_0872_ ), .B2(\myexu/myalu/_0396_ ), .ZN(\myexu/myalu/_0063_ ) );
AND3_X1 \myexu/myalu/_2349_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0385_ ), .ZN(\myexu/myalu/_0064_ ) );
OR4_X1 \myexu/myalu/_2350_ ( .A1(\myexu/myalu/_0044_ ), .A2(\myexu/myalu/_0061_ ), .A3(\myexu/myalu/_0063_ ), .A4(\myexu/myalu/_0064_ ), .ZN(\myexu/myalu/_1304_ ) );
AND2_X1 \myexu/myalu/_2351_ ( .A1(\myexu/myalu/_1062_ ), .A2(\myexu/myalu/_1063_ ), .ZN(\myexu/myalu/_0065_ ) );
AND2_X1 \myexu/myalu/_2352_ ( .A1(\myexu/myalu/_0864_ ), .A2(\myexu/myalu/_0865_ ), .ZN(\myexu/myalu/_0067_ ) );
OR2_X2 \myexu/myalu/_2353_ ( .A1(\myexu/myalu/_0065_ ), .A2(\myexu/myalu/_0067_ ), .ZN(\myexu/myalu/_0068_ ) );
INV_X1 \myexu/myalu/_2354_ ( .A(\myexu/myalu/_0046_ ), .ZN(\myexu/myalu/_0069_ ) );
NOR4_X1 \myexu/myalu/_2355_ ( .A1(\myexu/myalu/_0806_ ), .A2(\myexu/myalu/_0659_ ), .A3(\myexu/myalu/_0807_ ), .A4(\myexu/myalu/_0069_ ), .ZN(\myexu/myalu/_0070_ ) );
OAI21_X1 \myexu/myalu/_2356_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_0068_ ), .B2(\myexu/myalu/_0070_ ), .ZN(\myexu/myalu/_0071_ ) );
INV_X1 \myexu/myalu/_2357_ ( .A(\myexu/myalu/_0884_ ), .ZN(\myexu/myalu/_0072_ ) );
AOI21_X1 \myexu/myalu/_2358_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0072_ ), .B2(\myexu/myalu/_1386_ ), .ZN(\myexu/myalu/_0073_ ) );
NAND2_X1 \myexu/myalu/_2359_ ( .A1(\myexu/myalu/_1164_ ), .A2(\myexu/myalu/_1167_ ), .ZN(\myexu/myalu/_0074_ ) );
AOI21_X1 \myexu/myalu/_2360_ ( .A(\myexu/myalu/_0843_ ), .B1(\myexu/myalu/_1271_ ), .B2(\myexu/myalu/_1272_ ), .ZN(\myexu/myalu/_0075_ ) );
OR3_X1 \myexu/myalu/_2361_ ( .A1(\myexu/myalu/_0696_ ), .A2(\myexu/myalu/_0649_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_0076_ ) );
OR3_X1 \myexu/myalu/_2362_ ( .A1(\myexu/myalu/_0699_ ), .A2(\myexu/myalu/_0697_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0078_ ) );
AOI21_X1 \myexu/myalu/_2363_ ( .A(fanout_net_14 ), .B1(\myexu/myalu/_0076_ ), .B2(\myexu/myalu/_0078_ ), .ZN(\myexu/myalu/_0079_ ) );
NOR2_X1 \myexu/myalu/_2364_ ( .A1(\myexu/myalu/_0075_ ), .A2(\myexu/myalu/_0079_ ), .ZN(\myexu/myalu/_0080_ ) );
MUX2_X1 \myexu/myalu/_2365_ ( .A(\myexu/myalu/_0074_ ), .B(\myexu/myalu/_0080_ ), .S(\myexu/myalu/_0883_ ), .Z(\myexu/myalu/_0081_ ) );
OAI21_X1 \myexu/myalu/_2366_ ( .A(\myexu/myalu/_0073_ ), .B1(\myexu/myalu/_0081_ ), .B2(\myexu/myalu/_1386_ ), .ZN(\myexu/myalu/_0082_ ) );
NAND3_X1 \myexu/myalu/_2367_ ( .A1(\myexu/myalu/_0864_ ), .A2(\myexu/myalu/_0911_ ), .A3(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0083_ ) );
AND3_X1 \myexu/myalu/_2368_ ( .A1(\myexu/myalu/_0071_ ), .A2(\myexu/myalu/_0082_ ), .A3(\myexu/myalu/_0083_ ), .ZN(\myexu/myalu/_0084_ ) );
INV_X1 \myexu/myalu/_2369_ ( .A(\myexu/myalu/_0039_ ), .ZN(\myexu/myalu/_0085_ ) );
AOI21_X1 \myexu/myalu/_2370_ ( .A(\myexu/myalu/_0396_ ), .B1(\myexu/myalu/_0019_ ), .B2(\myexu/myalu/_0085_ ), .ZN(\myexu/myalu/_0086_ ) );
OR3_X1 \myexu/myalu/_2371_ ( .A1(\myexu/myalu/_0086_ ), .A2(\myexu/myalu/_0322_ ), .A3(\myexu/myalu/_0385_ ), .ZN(\myexu/myalu/_0087_ ) );
OAI21_X1 \myexu/myalu/_2372_ ( .A(\myexu/myalu/_0322_ ), .B1(\myexu/myalu/_0086_ ), .B2(\myexu/myalu/_0385_ ), .ZN(\myexu/myalu/_0089_ ) );
NAND3_X1 \myexu/myalu/_2373_ ( .A1(\myexu/myalu/_0087_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_0089_ ), .ZN(\myexu/myalu/_0090_ ) );
AOI21_X1 \myexu/myalu/_2374_ ( .A(\myexu/myalu/_0872_ ), .B1(\myexu/myalu/_0609_ ), .B2(\myexu/myalu/_0542_ ), .ZN(\myexu/myalu/_0091_ ) );
AOI21_X1 \myexu/myalu/_2375_ ( .A(\myexu/myalu/_0091_ ), .B1(\myexu/myalu/_0322_ ), .B2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_0092_ ) );
AND2_X1 \myexu/myalu/_2376_ ( .A1(\myexu/myalu/_1369_ ), .A2(\myexu/myalu/_1337_ ), .ZN(\myexu/myalu/_0093_ ) );
NAND3_X1 \myexu/myalu/_2377_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0093_ ), .ZN(\myexu/myalu/_0094_ ) );
NAND4_X1 \myexu/myalu/_2378_ ( .A1(\myexu/myalu/_0084_ ), .A2(\myexu/myalu/_0090_ ), .A3(\myexu/myalu/_0092_ ), .A4(\myexu/myalu/_0094_ ), .ZN(\myexu/myalu/_1305_ ) );
NAND2_X1 \myexu/myalu/_2379_ ( .A1(\myexu/myalu/_0908_ ), .A2(\myexu/myalu/_0911_ ), .ZN(\myexu/myalu/_0095_ ) );
OAI21_X1 \myexu/myalu/_2380_ ( .A(\myexu/myalu/_0095_ ), .B1(\myexu/myalu/_1260_ ), .B2(\myexu/myalu/_1261_ ), .ZN(\myexu/myalu/_0096_ ) );
NOR3_X1 \myexu/myalu/_2381_ ( .A1(\myexu/myalu/_0806_ ), .A2(\myexu/myalu/_0807_ ), .A3(\myexu/myalu/_0069_ ), .ZN(\myexu/myalu/_0097_ ) );
OAI21_X1 \myexu/myalu/_2382_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_0096_ ), .B2(\myexu/myalu/_0097_ ), .ZN(\myexu/myalu/_0099_ ) );
INV_X1 \myexu/myalu/_2383_ ( .A(\myexu/myalu/_0089_ ), .ZN(\myexu/myalu/_0100_ ) );
OR3_X1 \myexu/myalu/_2384_ ( .A1(\myexu/myalu/_0100_ ), .A2(\myexu/myalu/_0354_ ), .A3(\myexu/myalu/_0093_ ), .ZN(\myexu/myalu/_0101_ ) );
OAI21_X1 \myexu/myalu/_2385_ ( .A(\myexu/myalu/_0354_ ), .B1(\myexu/myalu/_0100_ ), .B2(\myexu/myalu/_0093_ ), .ZN(\myexu/myalu/_0102_ ) );
NAND3_X1 \myexu/myalu/_2386_ ( .A1(\myexu/myalu/_0101_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_0102_ ), .ZN(\myexu/myalu/_0103_ ) );
NOR4_X1 \myexu/myalu/_2387_ ( .A1(\myexu/myalu/_0343_ ), .A2(\myexu/myalu/_0675_ ), .A3(\myexu/myalu/_0000_ ), .A4(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0104_ ) );
AND3_X1 \myexu/myalu/_2388_ ( .A1(\myexu/myalu/_0908_ ), .A2(\myexu/myalu/_0866_ ), .A3(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_0105_ ) );
AOI211_X4 \myexu/myalu/_2389_ ( .A(\myexu/myalu/_0104_ ), .B(\myexu/myalu/_0105_ ), .C1(\myexu/myalu/_0354_ ), .C2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0106_ ) );
OR2_X1 \myexu/myalu/_2390_ ( .A1(\myexu/myalu/_0941_ ), .A2(fanout_net_16 ), .ZN(\myexu/myalu/_0107_ ) );
AOI21_X1 \myexu/myalu/_2391_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0107_ ), .B2(\myexu/myalu/_1386_ ), .ZN(\myexu/myalu/_0108_ ) );
AOI21_X1 \myexu/myalu/_2392_ ( .A(\myexu/myalu/_0873_ ), .B1(\myexu/myalu/_1288_ ), .B2(\myexu/myalu/_1289_ ), .ZN(\myexu/myalu/_0110_ ) );
OAI21_X1 \myexu/myalu/_2393_ ( .A(\myexu/myalu/_0839_ ), .B1(\myexu/myalu/_0735_ ), .B2(\myexu/myalu/_0739_ ), .ZN(\myexu/myalu/_0111_ ) );
OAI21_X1 \myexu/myalu/_2394_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0738_ ), .B2(\myexu/myalu/_0776_ ), .ZN(\myexu/myalu/_0112_ ) );
AND3_X1 \myexu/myalu/_2395_ ( .A1(\myexu/myalu/_0111_ ), .A2(\myexu/myalu/_0996_ ), .A3(\myexu/myalu/_0112_ ), .ZN(\myexu/myalu/_0113_ ) );
NOR3_X1 \myexu/myalu/_2396_ ( .A1(\myexu/myalu/_0110_ ), .A2(\myexu/myalu/_0113_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_0114_ ) );
AOI21_X1 \myexu/myalu/_2397_ ( .A(\myexu/myalu/_1000_ ), .B1(\myexu/myalu/_1187_ ), .B2(\myexu/myalu/_1190_ ), .ZN(\myexu/myalu/_0115_ ) );
OR3_X1 \myexu/myalu/_2398_ ( .A1(\myexu/myalu/_0114_ ), .A2(\myexu/myalu/_0115_ ), .A3(\myexu/myalu/_1386_ ), .ZN(\myexu/myalu/_0116_ ) );
AND2_X1 \myexu/myalu/_2399_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0729_ ), .ZN(\myexu/myalu/_0117_ ) );
AOI22_X1 \myexu/myalu/_2400_ ( .A1(\myexu/myalu/_0108_ ), .A2(\myexu/myalu/_0116_ ), .B1(\myexu/myalu/_0333_ ), .B2(\myexu/myalu/_0117_ ), .ZN(\myexu/myalu/_0118_ ) );
NAND4_X1 \myexu/myalu/_2401_ ( .A1(\myexu/myalu/_0099_ ), .A2(\myexu/myalu/_0103_ ), .A3(\myexu/myalu/_0106_ ), .A4(\myexu/myalu/_0118_ ), .ZN(\myexu/myalu/_1306_ ) );
AND2_X1 \myexu/myalu/_2402_ ( .A1(\myexu/myalu/_0417_ ), .A2(\myexu/myalu/_0407_ ), .ZN(\myexu/myalu/_0120_ ) );
AND3_X1 \myexu/myalu/_2403_ ( .A1(\myexu/myalu/_0120_ ), .A2(\myexu/myalu/_0354_ ), .A3(\myexu/myalu/_0322_ ), .ZN(\myexu/myalu/_0121_ ) );
INV_X1 \myexu/myalu/_2404_ ( .A(\myexu/myalu/_0121_ ), .ZN(\myexu/myalu/_0122_ ) );
AOI21_X2 \myexu/myalu/_2405_ ( .A(\myexu/myalu/_0122_ ), .B1(\myexu/myalu/_0012_ ), .B2(\myexu/myalu/_0017_ ), .ZN(\myexu/myalu/_0123_ ) );
NOR3_X1 \myexu/myalu/_2406_ ( .A1(\myexu/myalu/_0085_ ), .A2(\myexu/myalu/_0385_ ), .A3(\myexu/myalu/_0396_ ), .ZN(\myexu/myalu/_0124_ ) );
OAI211_X2 \myexu/myalu/_2407_ ( .A(\myexu/myalu/_0354_ ), .B(\myexu/myalu/_0322_ ), .C1(\myexu/myalu/_0124_ ), .C2(\myexu/myalu/_0385_ ), .ZN(\myexu/myalu/_0125_ ) );
AOI21_X1 \myexu/myalu/_2408_ ( .A(\myexu/myalu/_0333_ ), .B1(\myexu/myalu/_0354_ ), .B2(\myexu/myalu/_0093_ ), .ZN(\myexu/myalu/_0126_ ) );
AND2_X1 \myexu/myalu/_2409_ ( .A1(\myexu/myalu/_0125_ ), .A2(\myexu/myalu/_0126_ ), .ZN(\myexu/myalu/_0127_ ) );
INV_X1 \myexu/myalu/_2410_ ( .A(\myexu/myalu/_0127_ ), .ZN(\myexu/myalu/_0128_ ) );
OR3_X1 \myexu/myalu/_2411_ ( .A1(\myexu/myalu/_0123_ ), .A2(\myexu/myalu/_0268_ ), .A3(\myexu/myalu/_0128_ ), .ZN(\myexu/myalu/_0129_ ) );
OAI21_X1 \myexu/myalu/_2412_ ( .A(\myexu/myalu/_0268_ ), .B1(\myexu/myalu/_0123_ ), .B2(\myexu/myalu/_0128_ ), .ZN(\myexu/myalu/_0131_ ) );
AND3_X1 \myexu/myalu/_2413_ ( .A1(\myexu/myalu/_0129_ ), .A2(\myexu/myalu/_0827_ ), .A3(\myexu/myalu/_0131_ ), .ZN(\myexu/myalu/_0132_ ) );
NAND3_X1 \myexu/myalu/_2414_ ( .A1(\myexu/myalu/_0956_ ), .A2(\myexu/myalu/_0867_ ), .A3(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_0133_ ) );
AND4_X1 \myexu/myalu/_2415_ ( .A1(\myexu/myalu/_0633_ ), .A2(\myexu/myalu/_0803_ ), .A3(\myexu/myalu/_0805_ ), .A4(\myexu/myalu/_0046_ ), .ZN(\myexu/myalu/_0134_ ) );
AOI221_X1 \myexu/myalu/_2416_ ( .A(\myexu/myalu/_0134_ ), .B1(\myexu/myalu/_0865_ ), .B2(\myexu/myalu/_0956_ ), .C1(\myexu/myalu/_1062_ ), .C2(\myexu/myalu/_1063_ ), .ZN(\myexu/myalu/_0135_ ) );
OAI21_X1 \myexu/myalu/_2417_ ( .A(\myexu/myalu/_0133_ ), .B1(\myexu/myalu/_0135_ ), .B2(\myexu/myalu/_0950_ ), .ZN(\myexu/myalu/_0136_ ) );
NAND2_X1 \myexu/myalu/_2418_ ( .A1(\myexu/myalu/_0268_ ), .A2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0137_ ) );
OAI211_X2 \myexu/myalu/_2419_ ( .A(\myexu/myalu/_0676_ ), .B(\myexu/myalu/_0983_ ), .C1(\myexu/myalu/_1372_ ), .C2(\myexu/myalu/_1340_ ), .ZN(\myexu/myalu/_0138_ ) );
AND2_X1 \myexu/myalu/_2420_ ( .A1(\myexu/myalu/_1372_ ), .A2(\myexu/myalu/_1340_ ), .ZN(\myexu/myalu/_0139_ ) );
NAND3_X1 \myexu/myalu/_2421_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0983_ ), .A3(\myexu/myalu/_0139_ ), .ZN(\myexu/myalu/_0140_ ) );
NAND3_X1 \myexu/myalu/_2422_ ( .A1(\myexu/myalu/_0137_ ), .A2(\myexu/myalu/_0138_ ), .A3(\myexu/myalu/_0140_ ), .ZN(\myexu/myalu/_0142_ ) );
OAI21_X1 \myexu/myalu/_2423_ ( .A(fanout_net_16 ), .B1(\myexu/myalu/_1223_ ), .B2(\myexu/myalu/_1224_ ), .ZN(\myexu/myalu/_0143_ ) );
OR3_X1 \myexu/myalu/_2424_ ( .A1(\myexu/myalu/_0699_ ), .A2(\myexu/myalu/_0697_ ), .A3(\myexu/myalu/_0695_ ), .ZN(\myexu/myalu/_0144_ ) );
OR3_X1 \myexu/myalu/_2425_ ( .A1(\myexu/myalu/_0705_ ), .A2(\myexu/myalu/_0700_ ), .A3(fanout_net_12 ), .ZN(\myexu/myalu/_0145_ ) );
NAND3_X1 \myexu/myalu/_2426_ ( .A1(\myexu/myalu/_0144_ ), .A2(\myexu/myalu/_0145_ ), .A3(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_0146_ ) );
NAND3_X1 \myexu/myalu/_2427_ ( .A1(\myexu/myalu/_0027_ ), .A2(\myexu/myalu/_0028_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_0147_ ) );
NAND2_X1 \myexu/myalu/_2428_ ( .A1(\myexu/myalu/_0146_ ), .A2(\myexu/myalu/_0147_ ), .ZN(\myexu/myalu/_0148_ ) );
OAI211_X2 \myexu/myalu/_2429_ ( .A(\myexu/myalu/_0143_ ), .B(\myexu/myalu/_0910_ ), .C1(fanout_net_16 ), .C2(\myexu/myalu/_0148_ ), .ZN(\myexu/myalu/_0149_ ) );
NAND3_X1 \myexu/myalu/_2430_ ( .A1(\myexu/myalu/_0979_ ), .A2(\myexu/myalu/_1386_ ), .A3(\myexu/myalu/_0980_ ), .ZN(\myexu/myalu/_0150_ ) );
AOI21_X1 \myexu/myalu/_2431_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0149_ ), .B2(\myexu/myalu/_0150_ ), .ZN(\myexu/myalu/_0151_ ) );
OR4_X1 \myexu/myalu/_2432_ ( .A1(\myexu/myalu/_0132_ ), .A2(\myexu/myalu/_0136_ ), .A3(\myexu/myalu/_0142_ ), .A4(\myexu/myalu/_0151_ ), .ZN(\myexu/myalu/_1308_ ) );
NOR4_X1 \myexu/myalu/_2433_ ( .A1(\myexu/myalu/_0290_ ), .A2(\myexu/myalu/_0675_ ), .A3(\myexu/myalu/_0000_ ), .A4(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0153_ ) );
AND3_X1 \myexu/myalu/_2434_ ( .A1(\myexu/myalu/_0992_ ), .A2(\myexu/myalu/_0866_ ), .A3(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_0154_ ) );
AOI211_X4 \myexu/myalu/_2435_ ( .A(\myexu/myalu/_0153_ ), .B(\myexu/myalu/_0154_ ), .C1(\myexu/myalu/_0301_ ), .C2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0155_ ) );
INV_X1 \myexu/myalu/_2436_ ( .A(\myexu/myalu/_0139_ ), .ZN(\myexu/myalu/_0156_ ) );
AND3_X1 \myexu/myalu/_2437_ ( .A1(\myexu/myalu/_0131_ ), .A2(\myexu/myalu/_0301_ ), .A3(\myexu/myalu/_0156_ ), .ZN(\myexu/myalu/_0157_ ) );
AOI21_X1 \myexu/myalu/_2438_ ( .A(\myexu/myalu/_0301_ ), .B1(\myexu/myalu/_0131_ ), .B2(\myexu/myalu/_0156_ ), .ZN(\myexu/myalu/_0158_ ) );
OAI21_X1 \myexu/myalu/_2439_ ( .A(\myexu/myalu/_0827_ ), .B1(\myexu/myalu/_0157_ ), .B2(\myexu/myalu/_0158_ ), .ZN(\myexu/myalu/_0159_ ) );
NAND3_X1 \myexu/myalu/_2440_ ( .A1(\myexu/myalu/_1243_ ), .A2(fanout_net_16 ), .A3(\myexu/myalu/_1244_ ), .ZN(\myexu/myalu/_0160_ ) );
AND3_X1 \myexu/myalu/_2441_ ( .A1(\myexu/myalu/_0052_ ), .A2(fanout_net_14 ), .A3(\myexu/myalu/_0053_ ), .ZN(\myexu/myalu/_0161_ ) );
OAI21_X1 \myexu/myalu/_2442_ ( .A(fanout_net_12 ), .B1(\myexu/myalu/_0735_ ), .B2(\myexu/myalu/_0739_ ), .ZN(\myexu/myalu/_0163_ ) );
OAI21_X1 \myexu/myalu/_2443_ ( .A(\myexu/myalu/_0905_ ), .B1(\myexu/myalu/_0746_ ), .B2(\myexu/myalu/_0736_ ), .ZN(\myexu/myalu/_0164_ ) );
AOI21_X1 \myexu/myalu/_2444_ ( .A(fanout_net_14 ), .B1(\myexu/myalu/_0163_ ), .B2(\myexu/myalu/_0164_ ), .ZN(\myexu/myalu/_0165_ ) );
OR2_X1 \myexu/myalu/_2445_ ( .A1(\myexu/myalu/_0161_ ), .A2(\myexu/myalu/_0165_ ), .ZN(\myexu/myalu/_0166_ ) );
OAI211_X2 \myexu/myalu/_2446_ ( .A(\myexu/myalu/_0160_ ), .B(\myexu/myalu/_0866_ ), .C1(\myexu/myalu/_0166_ ), .C2(fanout_net_16 ), .ZN(\myexu/myalu/_0167_ ) );
NAND3_X1 \myexu/myalu/_2447_ ( .A1(\myexu/myalu/_1014_ ), .A2(\myexu/myalu/_1386_ ), .A3(\myexu/myalu/_0883_ ), .ZN(\myexu/myalu/_0168_ ) );
AOI21_X1 \myexu/myalu/_2448_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0167_ ), .B2(\myexu/myalu/_0168_ ), .ZN(\myexu/myalu/_0169_ ) );
AOI21_X1 \myexu/myalu/_2449_ ( .A(\myexu/myalu/_0169_ ), .B1(\myexu/myalu/_0279_ ), .B2(\myexu/myalu/_0117_ ), .ZN(\myexu/myalu/_0170_ ) );
AND2_X1 \myexu/myalu/_2450_ ( .A1(\myexu/myalu/_0159_ ), .A2(\myexu/myalu/_0170_ ), .ZN(\myexu/myalu/_0171_ ) );
AND4_X1 \myexu/myalu/_2451_ ( .A1(\myexu/myalu/_0634_ ), .A2(\myexu/myalu/_0803_ ), .A3(\myexu/myalu/_1003_ ), .A4(\myexu/myalu/_0046_ ), .ZN(\myexu/myalu/_0172_ ) );
AOI221_X4 \myexu/myalu/_2452_ ( .A(\myexu/myalu/_0172_ ), .B1(\myexu/myalu/_0867_ ), .B2(\myexu/myalu/_0992_ ), .C1(\myexu/myalu/_1062_ ), .C2(\myexu/myalu/_1063_ ), .ZN(\myexu/myalu/_0174_ ) );
OAI211_X2 \myexu/myalu/_2453_ ( .A(\myexu/myalu/_0155_ ), .B(\myexu/myalu/_0171_ ), .C1(\myexu/myalu/_0174_ ), .C2(\myexu/myalu/_0950_ ), .ZN(\myexu/myalu/_1309_ ) );
OAI211_X2 \myexu/myalu/_2454_ ( .A(\myexu/myalu/_1035_ ), .B(\myexu/myalu/_0046_ ), .C1(fanout_net_14 ), .C2(\myexu/myalu/_0660_ ), .ZN(\myexu/myalu/_0175_ ) );
AOI22_X1 \myexu/myalu/_2455_ ( .A1(\myexu/myalu/_1062_ ), .A2(\myexu/myalu/_1063_ ), .B1(\myexu/myalu/_0867_ ), .B2(\myexu/myalu/_1025_ ), .ZN(\myexu/myalu/_0176_ ) );
AOI21_X1 \myexu/myalu/_2456_ ( .A(\myexu/myalu/_0950_ ), .B1(\myexu/myalu/_0175_ ), .B2(\myexu/myalu/_0176_ ), .ZN(\myexu/myalu/_0177_ ) );
NAND3_X1 \myexu/myalu/_2457_ ( .A1(\myexu/myalu/_1047_ ), .A2(\myexu/myalu/_1386_ ), .A3(\myexu/myalu/_1091_ ), .ZN(\myexu/myalu/_0178_ ) );
NAND3_X1 \myexu/myalu/_2458_ ( .A1(\myexu/myalu/_1273_ ), .A2(\myexu/myalu/_1274_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_0179_ ) );
OR3_X1 \myexu/myalu/_2459_ ( .A1(\myexu/myalu/_0705_ ), .A2(\myexu/myalu/_0700_ ), .A3(\myexu/myalu/_0905_ ), .ZN(\myexu/myalu/_0180_ ) );
OR3_X1 \myexu/myalu/_2460_ ( .A1(\myexu/myalu/_0708_ ), .A2(\myexu/myalu/_0706_ ), .A3(\myexu/myalu/_1371_ ), .ZN(\myexu/myalu/_0181_ ) );
NAND3_X1 \myexu/myalu/_2461_ ( .A1(\myexu/myalu/_0180_ ), .A2(\myexu/myalu/_0181_ ), .A3(\myexu/myalu/_0843_ ), .ZN(\myexu/myalu/_0182_ ) );
NAND3_X1 \myexu/myalu/_2462_ ( .A1(\myexu/myalu/_0076_ ), .A2(\myexu/myalu/_0078_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_0184_ ) );
NAND2_X1 \myexu/myalu/_2463_ ( .A1(\myexu/myalu/_0182_ ), .A2(\myexu/myalu/_0184_ ), .ZN(\myexu/myalu/_0185_ ) );
OAI211_X2 \myexu/myalu/_2464_ ( .A(\myexu/myalu/_0179_ ), .B(\myexu/myalu/_0867_ ), .C1(\myexu/myalu/_0185_ ), .C2(fanout_net_16 ), .ZN(\myexu/myalu/_0186_ ) );
AOI21_X1 \myexu/myalu/_2465_ ( .A(\myexu/myalu/_0801_ ), .B1(\myexu/myalu/_0178_ ), .B2(\myexu/myalu/_0186_ ), .ZN(\myexu/myalu/_0187_ ) );
AND3_X1 \myexu/myalu/_2466_ ( .A1(\myexu/myalu/_1025_ ), .A2(\myexu/myalu/_0911_ ), .A3(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0188_ ) );
NOR3_X1 \myexu/myalu/_2467_ ( .A1(\myexu/myalu/_0177_ ), .A2(\myexu/myalu/_0187_ ), .A3(\myexu/myalu/_0188_ ), .ZN(\myexu/myalu/_0189_ ) );
AOI21_X1 \myexu/myalu/_2468_ ( .A(\myexu/myalu/_0290_ ), .B1(\myexu/myalu/_0131_ ), .B2(\myexu/myalu/_0156_ ), .ZN(\myexu/myalu/_0190_ ) );
OR3_X1 \myexu/myalu/_2469_ ( .A1(\myexu/myalu/_0190_ ), .A2(\myexu/myalu/_0215_ ), .A3(\myexu/myalu/_0279_ ), .ZN(\myexu/myalu/_0191_ ) );
OAI21_X1 \myexu/myalu/_2470_ ( .A(\myexu/myalu/_0215_ ), .B1(\myexu/myalu/_0190_ ), .B2(\myexu/myalu/_0279_ ), .ZN(\myexu/myalu/_0192_ ) );
NAND3_X1 \myexu/myalu/_2471_ ( .A1(\myexu/myalu/_0191_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_0192_ ), .ZN(\myexu/myalu/_0193_ ) );
NAND2_X1 \myexu/myalu/_2472_ ( .A1(\myexu/myalu/_0215_ ), .A2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_0195_ ) );
OAI211_X2 \myexu/myalu/_2473_ ( .A(\myexu/myalu/_0676_ ), .B(\myexu/myalu/_0822_ ), .C1(\myexu/myalu/_1374_ ), .C2(\myexu/myalu/_1342_ ), .ZN(\myexu/myalu/_0196_ ) );
AND2_X1 \myexu/myalu/_2474_ ( .A1(\myexu/myalu/_0195_ ), .A2(\myexu/myalu/_0196_ ), .ZN(\myexu/myalu/_0197_ ) );
AND2_X1 \myexu/myalu/_2475_ ( .A1(\myexu/myalu/_1374_ ), .A2(\myexu/myalu/_1342_ ), .ZN(\myexu/myalu/_0198_ ) );
NAND3_X1 \myexu/myalu/_2476_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0198_ ), .ZN(\myexu/myalu/_0199_ ) );
NAND4_X1 \myexu/myalu/_2477_ ( .A1(\myexu/myalu/_0189_ ), .A2(\myexu/myalu/_0193_ ), .A3(\myexu/myalu/_0197_ ), .A4(\myexu/myalu/_0199_ ), .ZN(\myexu/myalu/_1310_ ) );
INV_X1 \myexu/myalu/_2478_ ( .A(\myexu/myalu/_0192_ ), .ZN(\myexu/myalu/_0200_ ) );
OR3_X1 \myexu/myalu/_2479_ ( .A1(\myexu/myalu/_0200_ ), .A2(\myexu/myalu/_0247_ ), .A3(\myexu/myalu/_0198_ ), .ZN(\myexu/myalu/_0201_ ) );
OAI21_X1 \myexu/myalu/_2480_ ( .A(\myexu/myalu/_0247_ ), .B1(\myexu/myalu/_0200_ ), .B2(\myexu/myalu/_0198_ ), .ZN(\myexu/myalu/_0202_ ) );
AND3_X1 \myexu/myalu/_2481_ ( .A1(\myexu/myalu/_0201_ ), .A2(\myexu/myalu/_0827_ ), .A3(\myexu/myalu/_0202_ ), .ZN(\myexu/myalu/_0203_ ) );
AOI21_X1 \myexu/myalu/_2482_ ( .A(\myexu/myalu/_0882_ ), .B1(\myexu/myalu/_0584_ ), .B2(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_0205_ ) );
OR3_X1 \myexu/myalu/_2483_ ( .A1(\myexu/myalu/_0587_ ), .A2(\myexu/myalu/_1386_ ), .A3(\myexu/myalu/_0205_ ), .ZN(\myexu/myalu/_0206_ ) );
NAND4_X1 \myexu/myalu/_2484_ ( .A1(\myexu/myalu/_0634_ ), .A2(\myexu/myalu/_0810_ ), .A3(\myexu/myalu/_0815_ ), .A4(\myexu/myalu/_0206_ ), .ZN(\myexu/myalu/_0207_ ) );
NAND2_X1 \myexu/myalu/_2485_ ( .A1(\myexu/myalu/_1069_ ), .A2(\myexu/myalu/_0911_ ), .ZN(\myexu/myalu/_0208_ ) );
AOI21_X1 \myexu/myalu/_2486_ ( .A(\myexu/myalu/_0678_ ), .B1(\myexu/myalu/_0207_ ), .B2(\myexu/myalu/_0208_ ), .ZN(\myexu/myalu/_0209_ ) );
NAND2_X1 \myexu/myalu/_2487_ ( .A1(\myexu/myalu/_1290_ ), .A2(\myexu/myalu/_1291_ ), .ZN(\myexu/myalu/_0210_ ) );
NAND2_X1 \myexu/myalu/_2488_ ( .A1(\myexu/myalu/_0210_ ), .A2(fanout_net_16 ), .ZN(\myexu/myalu/_0211_ ) );
OAI21_X1 \myexu/myalu/_2489_ ( .A(\myexu/myalu/_0839_ ), .B1(\myexu/myalu/_0743_ ), .B2(\myexu/myalu/_0747_ ), .ZN(\myexu/myalu/_0212_ ) );
OAI21_X1 \myexu/myalu/_2490_ ( .A(\myexu/myalu/_1371_ ), .B1(\myexu/myalu/_0746_ ), .B2(\myexu/myalu/_0736_ ), .ZN(\myexu/myalu/_0213_ ) );
AOI21_X1 \myexu/myalu/_2491_ ( .A(fanout_net_14 ), .B1(\myexu/myalu/_0212_ ), .B2(\myexu/myalu/_0213_ ), .ZN(\myexu/myalu/_0214_ ) );
AOI21_X1 \myexu/myalu/_2492_ ( .A(\myexu/myalu/_0880_ ), .B1(\myexu/myalu/_0111_ ), .B2(\myexu/myalu/_0112_ ), .ZN(\myexu/myalu/_0216_ ) );
OAI21_X1 \myexu/myalu/_2493_ ( .A(\myexu/myalu/_0883_ ), .B1(\myexu/myalu/_0214_ ), .B2(\myexu/myalu/_0216_ ), .ZN(\myexu/myalu/_0217_ ) );
AOI21_X1 \myexu/myalu/_2494_ ( .A(\myexu/myalu/_0942_ ), .B1(\myexu/myalu/_0211_ ), .B2(\myexu/myalu/_0217_ ), .ZN(\myexu/myalu/_0218_ ) );
AND2_X1 \myexu/myalu/_2495_ ( .A1(\myexu/myalu/_0717_ ), .A2(\myexu/myalu/_1386_ ), .ZN(\myexu/myalu/_0219_ ) );
BUF_X2 \myexu/myalu/_2496_ ( .A(\myexu/myalu/_0219_ ), .Z(\myexu/myalu/_0220_ ) );
AND3_X1 \myexu/myalu/_2497_ ( .A1(\myexu/myalu/_1083_ ), .A2(\myexu/myalu/_0883_ ), .A3(\myexu/myalu/_0220_ ), .ZN(\myexu/myalu/_0221_ ) );
AND3_X1 \myexu/myalu/_2498_ ( .A1(\myexu/myalu/_0728_ ), .A2(\myexu/myalu/_0729_ ), .A3(\myexu/myalu/_0226_ ), .ZN(\myexu/myalu/_0222_ ) );
NAND3_X1 \myexu/myalu/_2499_ ( .A1(\myexu/myalu/_0247_ ), .A2(\myexu/myalu/_0572_ ), .A3(\myexu/myalu/_0635_ ), .ZN(\myexu/myalu/_0223_ ) );
OAI21_X1 \myexu/myalu/_2500_ ( .A(\myexu/myalu/_0223_ ), .B1(\myexu/myalu/_0872_ ), .B2(\myexu/myalu/_0236_ ), .ZN(\myexu/myalu/_0224_ ) );
OR4_X1 \myexu/myalu/_2501_ ( .A1(\myexu/myalu/_0218_ ), .A2(\myexu/myalu/_0221_ ), .A3(\myexu/myalu/_0222_ ), .A4(\myexu/myalu/_0224_ ), .ZN(\myexu/myalu/_0225_ ) );
OR3_X1 \myexu/myalu/_2502_ ( .A1(\myexu/myalu/_0203_ ), .A2(\myexu/myalu/_0209_ ), .A3(\myexu/myalu/_0225_ ), .ZN(\myexu/myalu/_1311_ ) );
AND3_X1 \myexu/myalu/_2503_ ( .A1(\myexu/myalu/_0634_ ), .A2(\myexu/myalu/_1089_ ), .A3(\myexu/myalu/_0046_ ), .ZN(\myexu/myalu/_0227_ ) );
AND2_X1 \myexu/myalu/_2504_ ( .A1(\myexu/myalu/_0693_ ), .A2(\myexu/myalu/_0995_ ), .ZN(\myexu/myalu/_0228_ ) );
AND2_X1 \myexu/myalu/_2505_ ( .A1(\myexu/myalu/_0228_ ), .A2(\myexu/myalu/_0910_ ), .ZN(\myexu/myalu/_0229_ ) );
OR2_X1 \myexu/myalu/_2506_ ( .A1(\myexu/myalu/_0227_ ), .A2(\myexu/myalu/_0229_ ), .ZN(\myexu/myalu/_0230_ ) );
OAI21_X1 \myexu/myalu/_2507_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_0230_ ), .B2(\myexu/myalu/_0065_ ), .ZN(\myexu/myalu/_0231_ ) );
AND2_X1 \myexu/myalu/_2508_ ( .A1(\myexu/myalu/_0268_ ), .A2(\myexu/myalu/_0301_ ), .ZN(\myexu/myalu/_0232_ ) );
AND2_X1 \myexu/myalu/_2509_ ( .A1(\myexu/myalu/_0215_ ), .A2(\myexu/myalu/_0247_ ), .ZN(\myexu/myalu/_0233_ ) );
AND2_X1 \myexu/myalu/_2510_ ( .A1(\myexu/myalu/_0232_ ), .A2(\myexu/myalu/_0233_ ), .ZN(\myexu/myalu/_0234_ ) );
NAND2_X1 \myexu/myalu/_2511_ ( .A1(\myexu/myalu/_0123_ ), .A2(\myexu/myalu/_0234_ ), .ZN(\myexu/myalu/_0235_ ) );
AND2_X1 \myexu/myalu/_2512_ ( .A1(\myexu/myalu/_0128_ ), .A2(\myexu/myalu/_0234_ ), .ZN(\myexu/myalu/_0237_ ) );
INV_X1 \myexu/myalu/_2513_ ( .A(\myexu/myalu/_0279_ ), .ZN(\myexu/myalu/_0238_ ) );
AOI21_X1 \myexu/myalu/_2514_ ( .A(\myexu/myalu/_0290_ ), .B1(\myexu/myalu/_0238_ ), .B2(\myexu/myalu/_0156_ ), .ZN(\myexu/myalu/_0239_ ) );
AND3_X1 \myexu/myalu/_2515_ ( .A1(\myexu/myalu/_0239_ ), .A2(\myexu/myalu/_0247_ ), .A3(\myexu/myalu/_0215_ ), .ZN(\myexu/myalu/_0240_ ) );
AND2_X1 \myexu/myalu/_2516_ ( .A1(\myexu/myalu/_0247_ ), .A2(\myexu/myalu/_0198_ ), .ZN(\myexu/myalu/_0241_ ) );
NOR4_X1 \myexu/myalu/_2517_ ( .A1(\myexu/myalu/_0237_ ), .A2(\myexu/myalu/_0226_ ), .A3(\myexu/myalu/_0240_ ), .A4(\myexu/myalu/_0241_ ), .ZN(\myexu/myalu/_0242_ ) );
NAND2_X1 \myexu/myalu/_2518_ ( .A1(\myexu/myalu/_0235_ ), .A2(\myexu/myalu/_0242_ ), .ZN(\myexu/myalu/_0243_ ) );
AND2_X1 \myexu/myalu/_2519_ ( .A1(\myexu/myalu/_0243_ ), .A2(\myexu/myalu/_0035_ ), .ZN(\myexu/myalu/_0244_ ) );
OAI21_X1 \myexu/myalu/_2520_ ( .A(\myexu/myalu/_0827_ ), .B1(\myexu/myalu/_0243_ ), .B2(\myexu/myalu/_0035_ ), .ZN(\myexu/myalu/_0245_ ) );
OR2_X1 \myexu/myalu/_2521_ ( .A1(\myexu/myalu/_0244_ ), .A2(\myexu/myalu/_0245_ ), .ZN(\myexu/myalu/_0246_ ) );
AOI21_X1 \myexu/myalu/_2522_ ( .A(\myexu/myalu/_0872_ ), .B1(\myexu/myalu/_0561_ ), .B2(\myexu/myalu/_0682_ ), .ZN(\myexu/myalu/_0248_ ) );
AOI221_X4 \myexu/myalu/_2523_ ( .A(\myexu/myalu/_0248_ ), .B1(\myexu/myalu/_0035_ ), .B2(\myexu/myalu/_0721_ ), .C1(\myexu/myalu/_0229_ ), .C2(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_0249_ ) );
NAND3_X1 \myexu/myalu/_2524_ ( .A1(\myexu/myalu/_0144_ ), .A2(\myexu/myalu/_0145_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_0250_ ) );
OR3_X1 \myexu/myalu/_2525_ ( .A1(\myexu/myalu/_0708_ ), .A2(\myexu/myalu/_0706_ ), .A3(\myexu/myalu/_0788_ ), .ZN(\myexu/myalu/_0251_ ) );
OAI211_X2 \myexu/myalu/_2526_ ( .A(\myexu/myalu/_0855_ ), .B(\myexu/myalu/_0695_ ), .C1(\myexu/myalu/_1360_ ), .C2(\myexu/myalu/_0682_ ), .ZN(\myexu/myalu/_0252_ ) );
AND2_X1 \myexu/myalu/_2527_ ( .A1(\myexu/myalu/_0251_ ), .A2(\myexu/myalu/_0252_ ), .ZN(\myexu/myalu/_0253_ ) );
INV_X1 \myexu/myalu/_2528_ ( .A(\myexu/myalu/_0253_ ), .ZN(\myexu/myalu/_0254_ ) );
OAI211_X2 \myexu/myalu/_2529_ ( .A(\myexu/myalu/_0995_ ), .B(\myexu/myalu/_0250_ ), .C1(\myexu/myalu/_0254_ ), .C2(fanout_net_14 ), .ZN(\myexu/myalu/_0255_ ) );
NAND3_X1 \myexu/myalu/_2530_ ( .A1(\myexu/myalu/_0029_ ), .A2(\myexu/myalu/_0030_ ), .A3(fanout_net_16 ), .ZN(\myexu/myalu/_0256_ ) );
AND3_X1 \myexu/myalu/_2531_ ( .A1(\myexu/myalu/_0255_ ), .A2(\myexu/myalu/_0885_ ), .A3(\myexu/myalu/_0256_ ), .ZN(\myexu/myalu/_0257_ ) );
AND2_X1 \myexu/myalu/_2532_ ( .A1(\myexu/myalu/_1376_ ), .A2(\myexu/myalu/_1344_ ), .ZN(\myexu/myalu/_0259_ ) );
AOI221_X4 \myexu/myalu/_2533_ ( .A(\myexu/myalu/_0257_ ), .B1(\myexu/myalu/_0259_ ), .B2(\myexu/myalu/_0117_ ), .C1(\myexu/myalu/_1112_ ), .C2(\myexu/myalu/_0220_ ), .ZN(\myexu/myalu/_0260_ ) );
NAND4_X1 \myexu/myalu/_2534_ ( .A1(\myexu/myalu/_0231_ ), .A2(\myexu/myalu/_0246_ ), .A3(\myexu/myalu/_0249_ ), .A4(\myexu/myalu/_0260_ ), .ZN(\myexu/myalu/_1312_ ) );
AND2_X2 \myexu/myalu/_2535_ ( .A1(\myexu/myalu/_0606_ ), .A2(\myexu/myalu/_0607_ ), .ZN(\myexu/myalu/_0261_ ) );
AND2_X1 \myexu/myalu/_2536_ ( .A1(\myexu/myalu/_0261_ ), .A2(\myexu/myalu/_0613_ ), .ZN(\myexu/myalu/_0262_ ) );
INV_X1 \myexu/myalu/_2537_ ( .A(\myexu/myalu/_0262_ ), .ZN(\myexu/myalu/_0263_ ) );
NOR2_X2 \myexu/myalu/_2538_ ( .A1(\myexu/myalu/_0263_ ), .A2(\myexu/myalu/_0618_ ), .ZN(\myexu/myalu/_0264_ ) );
AND3_X4 \myexu/myalu/_2539_ ( .A1(\myexu/myalu/_0606_ ), .A2(\myexu/myalu/_0607_ ), .A3(\myexu/myalu/_0610_ ), .ZN(\myexu/myalu/_0265_ ) );
AND2_X4 \myexu/myalu/_2540_ ( .A1(\myexu/myalu/_0265_ ), .A2(\myexu/myalu/_0611_ ), .ZN(\myexu/myalu/_0266_ ) );
INV_X1 \myexu/myalu/_2541_ ( .A(\myexu/myalu/_0266_ ), .ZN(\myexu/myalu/_0267_ ) );
INV_X2 \myexu/myalu/_2542_ ( .A(\myexu/myalu/_0261_ ), .ZN(\myexu/myalu/_0269_ ) );
AND4_X1 \myexu/myalu/_2543_ ( .A1(\myexu/myalu/_1367_ ), .A2(\myexu/myalu/_0623_ ), .A3(\myexu/myalu/_1369_ ), .A4(\myexu/myalu/_1370_ ), .ZN(\myexu/myalu/_0270_ ) );
NAND3_X1 \myexu/myalu/_2544_ ( .A1(\myexu/myalu/_0269_ ), .A2(\myexu/myalu/_1368_ ), .A3(\myexu/myalu/_0270_ ), .ZN(\myexu/myalu/_0271_ ) );
NAND2_X1 \myexu/myalu/_2545_ ( .A1(\myexu/myalu/_0267_ ), .A2(\myexu/myalu/_0271_ ), .ZN(\myexu/myalu/_0272_ ) );
INV_X1 \myexu/myalu/_2546_ ( .A(\myexu/myalu/_0612_ ), .ZN(\myexu/myalu/_0273_ ) );
AND3_X1 \myexu/myalu/_2547_ ( .A1(\myexu/myalu/_1364_ ), .A2(\myexu/myalu/_1365_ ), .A3(\myexu/myalu/_1366_ ), .ZN(\myexu/myalu/_0274_ ) );
NAND3_X1 \myexu/myalu/_2548_ ( .A1(\myexu/myalu/_0601_ ), .A2(\myexu/myalu/_1363_ ), .A3(\myexu/myalu/_0274_ ), .ZN(\myexu/myalu/_0275_ ) );
AOI22_X2 \myexu/myalu/_2549_ ( .A1(\myexu/myalu/_0266_ ), .A2(\myexu/myalu/_0273_ ), .B1(\myexu/myalu/_0269_ ), .B2(\myexu/myalu/_0275_ ), .ZN(\myexu/myalu/_0276_ ) );
NAND2_X1 \myexu/myalu/_2550_ ( .A1(\myexu/myalu/_0272_ ), .A2(\myexu/myalu/_0276_ ), .ZN(\myexu/myalu/_0277_ ) );
AND2_X1 \myexu/myalu/_2551_ ( .A1(\myexu/myalu/_1376_ ), .A2(\myexu/myalu/_1379_ ), .ZN(\myexu/myalu/_0278_ ) );
NAND4_X1 \myexu/myalu/_2552_ ( .A1(\myexu/myalu/_0625_ ), .A2(\myexu/myalu/_1377_ ), .A3(\myexu/myalu/_1378_ ), .A4(\myexu/myalu/_0278_ ), .ZN(\myexu/myalu/_0280_ ) );
AOI211_X2 \myexu/myalu/_2553_ ( .A(\myexu/myalu/_0264_ ), .B(\myexu/myalu/_0277_ ), .C1(\myexu/myalu/_0263_ ), .C2(\myexu/myalu/_0280_ ), .ZN(\myexu/myalu/_0281_ ) );
AND2_X2 \myexu/myalu/_2554_ ( .A1(\myexu/myalu/_0281_ ), .A2(\myexu/myalu/_0605_ ), .ZN(\myexu/myalu/_0282_ ) );
AND2_X4 \myexu/myalu/_2555_ ( .A1(\myexu/myalu/_0282_ ), .A2(\myexu/myalu/_0810_ ), .ZN(\myexu/myalu/_0283_ ) );
INV_X2 \myexu/myalu/_2556_ ( .A(\myexu/myalu/_0283_ ), .ZN(\myexu/myalu/_0284_ ) );
AOI21_X1 \myexu/myalu/_2557_ ( .A(\myexu/myalu/_0284_ ), .B1(\myexu/myalu/_1261_ ), .B2(\myexu/myalu/_1130_ ), .ZN(\myexu/myalu/_0285_ ) );
INV_X1 \myexu/myalu/_2558_ ( .A(\myexu/myalu/_0285_ ), .ZN(\myexu/myalu/_0286_ ) );
AOI21_X1 \myexu/myalu/_2559_ ( .A(\myexu/myalu/_0286_ ), .B1(\myexu/myalu/_1261_ ), .B2(\myexu/myalu/_1145_ ), .ZN(\myexu/myalu/_0287_ ) );
INV_X1 \myexu/myalu/_2560_ ( .A(\myexu/myalu/_0287_ ), .ZN(\myexu/myalu/_0288_ ) );
AOI21_X1 \myexu/myalu/_2561_ ( .A(\myexu/myalu/_0288_ ), .B1(\myexu/myalu/_1261_ ), .B2(\myexu/myalu/_1134_ ), .ZN(\myexu/myalu/_0289_ ) );
AND2_X1 \myexu/myalu/_2562_ ( .A1(\myexu/myalu/_0763_ ), .A2(\myexu/myalu/_0995_ ), .ZN(\myexu/myalu/_0291_ ) );
AND2_X1 \myexu/myalu/_2563_ ( .A1(\myexu/myalu/_0291_ ), .A2(\myexu/myalu/_0910_ ), .ZN(\myexu/myalu/_0292_ ) );
OAI21_X1 \myexu/myalu/_2564_ ( .A(\myexu/myalu/_0815_ ), .B1(\myexu/myalu/_0289_ ), .B2(\myexu/myalu/_0292_ ), .ZN(\myexu/myalu/_0293_ ) );
NAND3_X1 \myexu/myalu/_2565_ ( .A1(\myexu/myalu/_1126_ ), .A2(\myexu/myalu/_1127_ ), .A3(\myexu/myalu/_0220_ ), .ZN(\myexu/myalu/_0294_ ) );
AND3_X1 \myexu/myalu/_2566_ ( .A1(\myexu/myalu/_0163_ ), .A2(fanout_net_14 ), .A3(\myexu/myalu/_0164_ ), .ZN(\myexu/myalu/_0295_ ) );
OR3_X1 \myexu/myalu/_2567_ ( .A1(\myexu/myalu/_0743_ ), .A2(\myexu/myalu/_0905_ ), .A3(\myexu/myalu/_0747_ ), .ZN(\myexu/myalu/_0296_ ) );
OR3_X1 \myexu/myalu/_2568_ ( .A1(\myexu/myalu/_0756_ ), .A2(\myexu/myalu/_1371_ ), .A3(\myexu/myalu/_0744_ ), .ZN(\myexu/myalu/_0297_ ) );
NAND2_X1 \myexu/myalu/_2569_ ( .A1(\myexu/myalu/_0296_ ), .A2(\myexu/myalu/_0297_ ), .ZN(\myexu/myalu/_0298_ ) );
AOI211_X4 \myexu/myalu/_2570_ ( .A(fanout_net_16 ), .B(\myexu/myalu/_0295_ ), .C1(\myexu/myalu/_0873_ ), .C2(\myexu/myalu/_0298_ ), .ZN(\myexu/myalu/_0299_ ) );
AOI21_X1 \myexu/myalu/_2571_ ( .A(\myexu/myalu/_1000_ ), .B1(\myexu/myalu/_0051_ ), .B2(\myexu/myalu/_0054_ ), .ZN(\myexu/myalu/_0300_ ) );
OAI21_X1 \myexu/myalu/_2572_ ( .A(\myexu/myalu/_0886_ ), .B1(\myexu/myalu/_0299_ ), .B2(\myexu/myalu/_0300_ ), .ZN(\myexu/myalu/_0302_ ) );
NAND3_X1 \myexu/myalu/_2573_ ( .A1(\myexu/myalu/_0291_ ), .A2(\myexu/myalu/_0911_ ), .A3(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0303_ ) );
AND4_X2 \myexu/myalu/_2574_ ( .A1(\myexu/myalu/_0293_ ), .A2(\myexu/myalu/_0294_ ), .A3(\myexu/myalu/_0302_ ), .A4(\myexu/myalu/_0303_ ), .ZN(\myexu/myalu/_0304_ ) );
OR3_X1 \myexu/myalu/_2575_ ( .A1(\myexu/myalu/_0244_ ), .A2(\myexu/myalu/_0024_ ), .A3(\myexu/myalu/_0259_ ), .ZN(\myexu/myalu/_0305_ ) );
OAI21_X1 \myexu/myalu/_2576_ ( .A(\myexu/myalu/_0024_ ), .B1(\myexu/myalu/_0244_ ), .B2(\myexu/myalu/_0259_ ), .ZN(\myexu/myalu/_0306_ ) );
NAND3_X1 \myexu/myalu/_2577_ ( .A1(\myexu/myalu/_0305_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_0306_ ), .ZN(\myexu/myalu/_0307_ ) );
NOR4_X1 \myexu/myalu/_2578_ ( .A1(\myexu/myalu/_0013_ ), .A2(\myexu/myalu/_0675_ ), .A3(\myexu/myalu/_0000_ ), .A4(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0308_ ) );
AOI21_X1 \myexu/myalu/_2579_ ( .A(\myexu/myalu/_0308_ ), .B1(\myexu/myalu/_0024_ ), .B2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_0309_ ) );
NAND3_X1 \myexu/myalu/_2580_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0003_ ), .ZN(\myexu/myalu/_0310_ ) );
NAND4_X1 \myexu/myalu/_2581_ ( .A1(\myexu/myalu/_0304_ ), .A2(\myexu/myalu/_0307_ ), .A3(\myexu/myalu/_0309_ ), .A4(\myexu/myalu/_0310_ ), .ZN(\myexu/myalu/_1313_ ) );
OAI21_X1 \myexu/myalu/_2582_ ( .A(\myexu/myalu/_1062_ ), .B1(\myexu/myalu/_1063_ ), .B2(\myexu/myalu/_1131_ ), .ZN(\myexu/myalu/_0312_ ) );
AOI21_X1 \myexu/myalu/_2583_ ( .A(\myexu/myalu/_0312_ ), .B1(\myexu/myalu/_1261_ ), .B2(\myexu/myalu/_1145_ ), .ZN(\myexu/myalu/_0313_ ) );
AND2_X1 \myexu/myalu/_2584_ ( .A1(\myexu/myalu/_0863_ ), .A2(\myexu/myalu/_0995_ ), .ZN(\myexu/myalu/_0314_ ) );
AND2_X1 \myexu/myalu/_2585_ ( .A1(\myexu/myalu/_0314_ ), .A2(\myexu/myalu/_0910_ ), .ZN(\myexu/myalu/_0315_ ) );
OAI21_X1 \myexu/myalu/_2586_ ( .A(\myexu/myalu/_0815_ ), .B1(\myexu/myalu/_0313_ ), .B2(\myexu/myalu/_0315_ ), .ZN(\myexu/myalu/_0316_ ) );
NAND3_X1 \myexu/myalu/_2587_ ( .A1(\myexu/myalu/_0314_ ), .A2(\myexu/myalu/_0867_ ), .A3(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0317_ ) );
OAI211_X2 \myexu/myalu/_2588_ ( .A(\myexu/myalu/_0676_ ), .B(\myexu/myalu/_0945_ ), .C1(\myexu/myalu/_1378_ ), .C2(\myexu/myalu/_1346_ ), .ZN(\myexu/myalu/_0318_ ) );
NAND2_X1 \myexu/myalu/_2589_ ( .A1(\myexu/myalu/_0045_ ), .A2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0319_ ) );
AND4_X2 \myexu/myalu/_2590_ ( .A1(\myexu/myalu/_0316_ ), .A2(\myexu/myalu/_0317_ ), .A3(\myexu/myalu/_0318_ ), .A4(\myexu/myalu/_0319_ ), .ZN(\myexu/myalu/_0320_ ) );
NAND3_X1 \myexu/myalu/_2591_ ( .A1(\myexu/myalu/_0180_ ), .A2(\myexu/myalu/_0181_ ), .A3(fanout_net_14 ), .ZN(\myexu/myalu/_0321_ ) );
NOR2_X1 \myexu/myalu/_2592_ ( .A1(\myexu/myalu/_0679_ ), .A2(\myexu/myalu/_0684_ ), .ZN(\myexu/myalu/_0323_ ) );
NOR2_X1 \myexu/myalu/_2593_ ( .A1(\myexu/myalu/_0683_ ), .A2(\myexu/myalu/_0709_ ), .ZN(\myexu/myalu/_0324_ ) );
MUX2_X1 \myexu/myalu/_2594_ ( .A(\myexu/myalu/_0323_ ), .B(\myexu/myalu/_0324_ ), .S(\myexu/myalu/_1371_ ), .Z(\myexu/myalu/_0325_ ) );
OAI211_X2 \myexu/myalu/_2595_ ( .A(\myexu/myalu/_0980_ ), .B(\myexu/myalu/_0321_ ), .C1(\myexu/myalu/_0325_ ), .C2(fanout_net_14 ), .ZN(\myexu/myalu/_0326_ ) );
OAI211_X2 \myexu/myalu/_2596_ ( .A(\myexu/myalu/_0326_ ), .B(\myexu/myalu/_0886_ ), .C1(\myexu/myalu/_0080_ ), .C2(\myexu/myalu/_1091_ ), .ZN(\myexu/myalu/_0327_ ) );
OAI211_X2 \myexu/myalu/_2597_ ( .A(\myexu/myalu/_1168_ ), .B(\myexu/myalu/_0220_ ), .C1(\myexu/myalu/_0881_ ), .C2(\myexu/myalu/_1091_ ), .ZN(\myexu/myalu/_0328_ ) );
AND2_X1 \myexu/myalu/_2598_ ( .A1(\myexu/myalu/_1378_ ), .A2(\myexu/myalu/_1346_ ), .ZN(\myexu/myalu/_0329_ ) );
NAND3_X1 \myexu/myalu/_2599_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0329_ ), .ZN(\myexu/myalu/_0330_ ) );
AND3_X1 \myexu/myalu/_2600_ ( .A1(\myexu/myalu/_0327_ ), .A2(\myexu/myalu/_0328_ ), .A3(\myexu/myalu/_0330_ ), .ZN(\myexu/myalu/_0331_ ) );
NAND3_X1 \myexu/myalu/_2601_ ( .A1(\myexu/myalu/_0243_ ), .A2(\myexu/myalu/_0024_ ), .A3(\myexu/myalu/_0035_ ), .ZN(\myexu/myalu/_0332_ ) );
AOI21_X1 \myexu/myalu/_2602_ ( .A(\myexu/myalu/_0003_ ), .B1(\myexu/myalu/_0024_ ), .B2(\myexu/myalu/_0259_ ), .ZN(\myexu/myalu/_0334_ ) );
AND2_X1 \myexu/myalu/_2603_ ( .A1(\myexu/myalu/_0332_ ), .A2(\myexu/myalu/_0334_ ), .ZN(\myexu/myalu/_0335_ ) );
INV_X1 \myexu/myalu/_2604_ ( .A(\myexu/myalu/_0335_ ), .ZN(\myexu/myalu/_0336_ ) );
AND2_X1 \myexu/myalu/_2605_ ( .A1(\myexu/myalu/_0336_ ), .A2(\myexu/myalu/_0045_ ), .ZN(\myexu/myalu/_0337_ ) );
OAI21_X1 \myexu/myalu/_2606_ ( .A(\myexu/myalu/_0828_ ), .B1(\myexu/myalu/_0336_ ), .B2(\myexu/myalu/_0045_ ), .ZN(\myexu/myalu/_0338_ ) );
OAI211_X2 \myexu/myalu/_2607_ ( .A(\myexu/myalu/_0320_ ), .B(\myexu/myalu/_0331_ ), .C1(\myexu/myalu/_0337_ ), .C2(\myexu/myalu/_0338_ ), .ZN(\myexu/myalu/_1314_ ) );
NAND2_X1 \myexu/myalu/_2608_ ( .A1(\myexu/myalu/_1181_ ), .A2(\myexu/myalu/_0910_ ), .ZN(\myexu/myalu/_0339_ ) );
AOI21_X1 \myexu/myalu/_2609_ ( .A(\myexu/myalu/_0950_ ), .B1(\myexu/myalu/_0312_ ), .B2(\myexu/myalu/_0339_ ), .ZN(\myexu/myalu/_0340_ ) );
AND3_X1 \myexu/myalu/_2610_ ( .A1(\myexu/myalu/_1181_ ), .A2(\myexu/myalu/_0910_ ), .A3(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_0341_ ) );
NOR2_X1 \myexu/myalu/_2611_ ( .A1(\myexu/myalu/_0340_ ), .A2(\myexu/myalu/_0341_ ), .ZN(\myexu/myalu/_0342_ ) );
NAND3_X1 \myexu/myalu/_2612_ ( .A1(\myexu/myalu/_1186_ ), .A2(\myexu/myalu/_1191_ ), .A3(\myexu/myalu/_0220_ ), .ZN(\myexu/myalu/_0344_ ) );
OAI21_X1 \myexu/myalu/_2613_ ( .A(\myexu/myalu/_1385_ ), .B1(\myexu/myalu/_0110_ ), .B2(\myexu/myalu/_0113_ ), .ZN(\myexu/myalu/_0345_ ) );
NAND2_X1 \myexu/myalu/_2614_ ( .A1(\myexu/myalu/_0212_ ), .A2(\myexu/myalu/_0213_ ), .ZN(\myexu/myalu/_0346_ ) );
OR3_X1 \myexu/myalu/_2615_ ( .A1(\myexu/myalu/_0756_ ), .A2(\myexu/myalu/_0788_ ), .A3(\myexu/myalu/_0744_ ), .ZN(\myexu/myalu/_0347_ ) );
OR3_X1 \myexu/myalu/_2616_ ( .A1(\myexu/myalu/_0759_ ), .A2(\myexu/myalu/_0757_ ), .A3(\myexu/myalu/_1371_ ), .ZN(\myexu/myalu/_0348_ ) );
AND2_X1 \myexu/myalu/_2617_ ( .A1(\myexu/myalu/_0347_ ), .A2(\myexu/myalu/_0348_ ), .ZN(\myexu/myalu/_0349_ ) );
MUX2_X1 \myexu/myalu/_2618_ ( .A(\myexu/myalu/_0346_ ), .B(\myexu/myalu/_0349_ ), .S(\myexu/myalu/_0873_ ), .Z(\myexu/myalu/_0350_ ) );
OAI211_X2 \myexu/myalu/_2619_ ( .A(\myexu/myalu/_0886_ ), .B(\myexu/myalu/_0345_ ), .C1(\myexu/myalu/_0350_ ), .C2(\myexu/myalu/_1385_ ), .ZN(\myexu/myalu/_0351_ ) );
AND3_X1 \myexu/myalu/_2620_ ( .A1(\myexu/myalu/_0342_ ), .A2(\myexu/myalu/_0344_ ), .A3(\myexu/myalu/_0351_ ), .ZN(\myexu/myalu/_0352_ ) );
OR3_X1 \myexu/myalu/_2621_ ( .A1(\myexu/myalu/_0337_ ), .A2(\myexu/myalu/_0077_ ), .A3(\myexu/myalu/_0329_ ), .ZN(\myexu/myalu/_0353_ ) );
OAI21_X1 \myexu/myalu/_2622_ ( .A(\myexu/myalu/_0077_ ), .B1(\myexu/myalu/_0337_ ), .B2(\myexu/myalu/_0329_ ), .ZN(\myexu/myalu/_0355_ ) );
NAND3_X1 \myexu/myalu/_2623_ ( .A1(\myexu/myalu/_0353_ ), .A2(\myexu/myalu/_0828_ ), .A3(\myexu/myalu/_0355_ ), .ZN(\myexu/myalu/_0356_ ) );
NAND3_X1 \myexu/myalu/_2624_ ( .A1(\myexu/myalu/_0821_ ), .A2(\myexu/myalu/_0822_ ), .A3(\myexu/myalu/_0056_ ), .ZN(\myexu/myalu/_0357_ ) );
NOR4_X1 \myexu/myalu/_2625_ ( .A1(\myexu/myalu/_0066_ ), .A2(\myexu/myalu/_0675_ ), .A3(\myexu/myalu/_0000_ ), .A4(\myexu/myalu/_0002_ ), .ZN(\myexu/myalu/_0358_ ) );
AOI21_X1 \myexu/myalu/_2626_ ( .A(\myexu/myalu/_0358_ ), .B1(\myexu/myalu/_0077_ ), .B2(\myexu/myalu/_0819_ ), .ZN(\myexu/myalu/_0359_ ) );
NAND4_X1 \myexu/myalu/_2627_ ( .A1(\myexu/myalu/_0352_ ), .A2(\myexu/myalu/_0356_ ), .A3(\myexu/myalu/_0357_ ), .A4(\myexu/myalu/_0359_ ), .ZN(\myexu/myalu/_1315_ ) );
AND3_X2 \myexu/myalu/_2628_ ( .A1(\myexu/myalu/_0336_ ), .A2(\myexu/myalu/_0077_ ), .A3(\myexu/myalu/_0045_ ), .ZN(\myexu/myalu/_0360_ ) );
INV_X1 \myexu/myalu/_2629_ ( .A(\myexu/myalu/_0360_ ), .ZN(\myexu/myalu/_0361_ ) );
AOI21_X1 \myexu/myalu/_2630_ ( .A(\myexu/myalu/_0056_ ), .B1(\myexu/myalu/_0077_ ), .B2(\myexu/myalu/_0329_ ), .ZN(\myexu/myalu/_0362_ ) );
AND2_X2 \myexu/myalu/_2631_ ( .A1(\myexu/myalu/_0361_ ), .A2(\myexu/myalu/_0362_ ), .ZN(\myexu/myalu/_0363_ ) );
AOI21_X1 \myexu/myalu/_2632_ ( .A(\myexu/myalu/_0932_ ), .B1(\myexu/myalu/_0363_ ), .B2(\myexu/myalu/_0183_ ), .ZN(\myexu/myalu/_0365_ ) );
OAI21_X1 \myexu/myalu/_2633_ ( .A(\myexu/myalu/_0365_ ), .B1(\myexu/myalu/_0183_ ), .B2(\myexu/myalu/_0363_ ), .ZN(\myexu/myalu/_0366_ ) );
AND3_X1 \myexu/myalu/_2634_ ( .A1(\myexu/myalu/_0692_ ), .A2(\myexu/myalu/_0995_ ), .A3(\myexu/myalu/_0996_ ), .ZN(\myexu/myalu/_0367_ ) );
AND2_X1 \myexu/myalu/_2635_ ( .A1(\myexu/myalu/_0367_ ), .A2(\myexu/myalu/_0910_ ), .ZN(\myexu/myalu/_0368_ ) );
OR2_X1 \myexu/myalu/_2636_ ( .A1(\myexu/myalu/_0065_ ), .A2(\myexu/myalu/_0368_ ), .ZN(\myexu/myalu/_0369_ ) );
OR3_X1 \myexu/myalu/_2637_ ( .A1(\myexu/myalu/_0621_ ), .A2(\myexu/myalu/_0632_ ), .A3(\myexu/myalu/_0069_ ), .ZN(\myexu/myalu/_0370_ ) );
AOI21_X1 \myexu/myalu/_2638_ ( .A(\myexu/myalu/_0370_ ), .B1(\myexu/myalu/_1091_ ), .B2(\myexu/myalu/_0804_ ), .ZN(\myexu/myalu/_0371_ ) );
OAI21_X1 \myexu/myalu/_2639_ ( .A(\myexu/myalu/_0830_ ), .B1(\myexu/myalu/_0369_ ), .B2(\myexu/myalu/_0371_ ), .ZN(\myexu/myalu/_0372_ ) );
NAND2_X1 \myexu/myalu/_2640_ ( .A1(\myexu/myalu/_1226_ ), .A2(\myexu/myalu/_0220_ ), .ZN(\myexu/myalu/_0373_ ) );
NOR2_X1 \myexu/myalu/_2641_ ( .A1(\myexu/myalu/_0689_ ), .A2(\myexu/myalu/_0680_ ), .ZN(\myexu/myalu/_0374_ ) );
MUX2_X1 \myexu/myalu/_2642_ ( .A(\myexu/myalu/_0374_ ), .B(\myexu/myalu/_0323_ ), .S(\myexu/myalu/_1371_ ), .Z(\myexu/myalu/_0376_ ) );
MUX2_X1 \myexu/myalu/_2643_ ( .A(\myexu/myalu/_0376_ ), .B(\myexu/myalu/_0254_ ), .S(fanout_net_14 ), .Z(\myexu/myalu/_0377_ ) );
AOI21_X1 \myexu/myalu/_2644_ ( .A(\myexu/myalu/_0942_ ), .B1(\myexu/myalu/_0377_ ), .B2(\myexu/myalu/_0980_ ), .ZN(\myexu/myalu/_0378_ ) );
OAI21_X1 \myexu/myalu/_2645_ ( .A(\myexu/myalu/_0378_ ), .B1(\myexu/myalu/_1091_ ), .B2(\myexu/myalu/_0148_ ), .ZN(\myexu/myalu/_0379_ ) );
OAI21_X1 \myexu/myalu/_2646_ ( .A(\myexu/myalu/_0817_ ), .B1(\myexu/myalu/_1380_ ), .B2(\myexu/myalu/_1348_ ), .ZN(\myexu/myalu/_0380_ ) );
AND2_X1 \myexu/myalu/_2647_ ( .A1(\myexu/myalu/_1380_ ), .A2(\myexu/myalu/_1348_ ), .ZN(\myexu/myalu/_0381_ ) );
AOI22_X1 \myexu/myalu/_2648_ ( .A1(\myexu/myalu/_0117_ ), .A2(\myexu/myalu/_0381_ ), .B1(\myexu/myalu/_0173_ ), .B2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0382_ ) );
NAND3_X1 \myexu/myalu/_2649_ ( .A1(\myexu/myalu/_0367_ ), .A2(\myexu/myalu/_0867_ ), .A3(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0383_ ) );
AND4_X1 \myexu/myalu/_2650_ ( .A1(\myexu/myalu/_0379_ ), .A2(\myexu/myalu/_0380_ ), .A3(\myexu/myalu/_0382_ ), .A4(\myexu/myalu/_0383_ ), .ZN(\myexu/myalu/_0384_ ) );
NAND4_X1 \myexu/myalu/_2651_ ( .A1(\myexu/myalu/_0366_ ), .A2(\myexu/myalu/_0372_ ), .A3(\myexu/myalu/_0373_ ), .A4(\myexu/myalu/_0384_ ), .ZN(\myexu/myalu/_1316_ ) );
OAI211_X2 \myexu/myalu/_2652_ ( .A(\myexu/myalu/_0633_ ), .B(\myexu/myalu/_0046_ ), .C1(\myexu/myalu/_0803_ ), .C2(\myexu/myalu/_1003_ ), .ZN(\myexu/myalu/_0386_ ) );
INV_X1 \myexu/myalu/_2653_ ( .A(\myexu/myalu/_0386_ ), .ZN(\myexu/myalu/_0387_ ) );
AND3_X1 \myexu/myalu/_2654_ ( .A1(\myexu/myalu/_0755_ ), .A2(\myexu/myalu/_0505_ ), .A3(\myexu/myalu/_0773_ ), .ZN(\myexu/myalu/_0388_ ) );
AOI221_X1 \myexu/myalu/_2655_ ( .A(\myexu/myalu/_0387_ ), .B1(\myexu/myalu/_0865_ ), .B2(\myexu/myalu/_0388_ ), .C1(\myexu/myalu/_1062_ ), .C2(\myexu/myalu/_0811_ ), .ZN(\myexu/myalu/_0389_ ) );
OR2_X1 \myexu/myalu/_2656_ ( .A1(\myexu/myalu/_0389_ ), .A2(\myexu/myalu/_0950_ ), .ZN(\myexu/myalu/_0390_ ) );
OAI21_X1 \myexu/myalu/_2657_ ( .A(\myexu/myalu/_0220_ ), .B1(\myexu/myalu/_1239_ ), .B2(\myexu/myalu/_1245_ ), .ZN(\myexu/myalu/_0391_ ) );
NAND3_X1 \myexu/myalu/_2658_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0130_ ), .ZN(\myexu/myalu/_0392_ ) );
AND3_X1 \myexu/myalu/_2659_ ( .A1(\myexu/myalu/_0388_ ), .A2(\myexu/myalu/_0588_ ), .A3(\myexu/myalu/_0677_ ), .ZN(\myexu/myalu/_0393_ ) );
INV_X1 \myexu/myalu/_2660_ ( .A(\myexu/myalu/_0141_ ), .ZN(\myexu/myalu/_0394_ ) );
AOI221_X4 \myexu/myalu/_2661_ ( .A(\myexu/myalu/_0393_ ), .B1(\myexu/myalu/_0394_ ), .B2(\myexu/myalu/_0726_ ), .C1(\myexu/myalu/_0152_ ), .C2(\myexu/myalu/_0721_ ), .ZN(\myexu/myalu/_0395_ ) );
AND4_X2 \myexu/myalu/_2662_ ( .A1(\myexu/myalu/_0390_ ), .A2(\myexu/myalu/_0391_ ), .A3(\myexu/myalu/_0392_ ), .A4(\myexu/myalu/_0395_ ), .ZN(\myexu/myalu/_0397_ ) );
OR3_X1 \myexu/myalu/_2663_ ( .A1(\myexu/myalu/_0759_ ), .A2(\myexu/myalu/_0757_ ), .A3(\myexu/myalu/_0839_ ), .ZN(\myexu/myalu/_0398_ ) );
MUX2_X1 \myexu/myalu/_2664_ ( .A(\myexu/myalu/_1349_ ), .B(\myexu/myalu/_1348_ ), .S(\myexu/myalu/_1360_ ), .Z(\myexu/myalu/_0399_ ) );
OAI211_X2 \myexu/myalu/_2665_ ( .A(\myexu/myalu/_0398_ ), .B(\myexu/myalu/_0873_ ), .C1(\myexu/myalu/_1371_ ), .C2(\myexu/myalu/_0399_ ), .ZN(\myexu/myalu/_0400_ ) );
OAI21_X1 \myexu/myalu/_2666_ ( .A(\myexu/myalu/_0400_ ), .B1(\myexu/myalu/_0298_ ), .B2(\myexu/myalu/_0873_ ), .ZN(\myexu/myalu/_0401_ ) );
MUX2_X1 \myexu/myalu/_2667_ ( .A(\myexu/myalu/_0401_ ), .B(\myexu/myalu/_0166_ ), .S(\myexu/myalu/_1385_ ), .Z(\myexu/myalu/_0402_ ) );
NAND2_X1 \myexu/myalu/_2668_ ( .A1(\myexu/myalu/_0402_ ), .A2(\myexu/myalu/_0886_ ), .ZN(\myexu/myalu/_0403_ ) );
NOR2_X2 \myexu/myalu/_2669_ ( .A1(\myexu/myalu/_0363_ ), .A2(\myexu/myalu/_0183_ ), .ZN(\myexu/myalu/_0404_ ) );
INV_X1 \myexu/myalu/_2670_ ( .A(\myexu/myalu/_0404_ ), .ZN(\myexu/myalu/_0405_ ) );
INV_X1 \myexu/myalu/_2671_ ( .A(\myexu/myalu/_0381_ ), .ZN(\myexu/myalu/_0406_ ) );
NAND3_X1 \myexu/myalu/_2672_ ( .A1(\myexu/myalu/_0405_ ), .A2(\myexu/myalu/_0162_ ), .A3(\myexu/myalu/_0406_ ), .ZN(\myexu/myalu/_0408_ ) );
NAND2_X1 \myexu/myalu/_2673_ ( .A1(\myexu/myalu/_0408_ ), .A2(\myexu/myalu/_0828_ ), .ZN(\myexu/myalu/_0409_ ) );
AOI21_X1 \myexu/myalu/_2674_ ( .A(\myexu/myalu/_0162_ ), .B1(\myexu/myalu/_0405_ ), .B2(\myexu/myalu/_0406_ ), .ZN(\myexu/myalu/_0410_ ) );
OAI211_X2 \myexu/myalu/_2675_ ( .A(\myexu/myalu/_0397_ ), .B(\myexu/myalu/_0403_ ), .C1(\myexu/myalu/_0409_ ), .C2(\myexu/myalu/_0410_ ), .ZN(\myexu/myalu/_1317_ ) );
OR3_X2 \myexu/myalu/_2676_ ( .A1(\myexu/myalu/_0404_ ), .A2(\myexu/myalu/_0130_ ), .A3(\myexu/myalu/_0381_ ), .ZN(\myexu/myalu/_0411_ ) );
AND3_X1 \myexu/myalu/_2677_ ( .A1(\myexu/myalu/_0411_ ), .A2(\myexu/myalu/_0109_ ), .A3(\myexu/myalu/_0394_ ), .ZN(\myexu/myalu/_0412_ ) );
AOI21_X1 \myexu/myalu/_2678_ ( .A(\myexu/myalu/_0109_ ), .B1(\myexu/myalu/_0411_ ), .B2(\myexu/myalu/_0394_ ), .ZN(\myexu/myalu/_0413_ ) );
OR3_X1 \myexu/myalu/_2679_ ( .A1(\myexu/myalu/_0412_ ), .A2(\myexu/myalu/_0413_ ), .A3(\myexu/myalu/_0932_ ), .ZN(\myexu/myalu/_0414_ ) );
OR4_X1 \myexu/myalu/_2680_ ( .A1(\myexu/myalu/_0632_ ), .A2(\myexu/myalu/_0621_ ), .A3(\myexu/myalu/_1262_ ), .A4(\myexu/myalu/_0069_ ), .ZN(\myexu/myalu/_0415_ ) );
AND2_X1 \myexu/myalu/_2681_ ( .A1(\myexu/myalu/_1021_ ), .A2(\myexu/myalu/_1000_ ), .ZN(\myexu/myalu/_0416_ ) );
NAND2_X1 \myexu/myalu/_2682_ ( .A1(\myexu/myalu/_0416_ ), .A2(\myexu/myalu/_0911_ ), .ZN(\myexu/myalu/_0418_ ) );
OAI211_X2 \myexu/myalu/_2683_ ( .A(\myexu/myalu/_0415_ ), .B(\myexu/myalu/_0418_ ), .C1(\myexu/myalu/_1260_ ), .C2(\myexu/myalu/_1261_ ), .ZN(\myexu/myalu/_0419_ ) );
NAND2_X1 \myexu/myalu/_2684_ ( .A1(\myexu/myalu/_0419_ ), .A2(\myexu/myalu/_0830_ ), .ZN(\myexu/myalu/_0420_ ) );
OAI21_X1 \myexu/myalu/_2685_ ( .A(\myexu/myalu/_0220_ ), .B1(\myexu/myalu/_1270_ ), .B2(\myexu/myalu/_1275_ ), .ZN(\myexu/myalu/_0421_ ) );
OR3_X1 \myexu/myalu/_2686_ ( .A1(\myexu/myalu/_0689_ ), .A2(\myexu/myalu/_0680_ ), .A3(\myexu/myalu/_0905_ ), .ZN(\myexu/myalu/_0422_ ) );
MUX2_X1 \myexu/myalu/_2687_ ( .A(\myexu/myalu/_1351_ ), .B(\myexu/myalu/_1349_ ), .S(\myexu/myalu/_1360_ ), .Z(\myexu/myalu/_0423_ ) );
OAI211_X2 \myexu/myalu/_2688_ ( .A(\myexu/myalu/_0422_ ), .B(\myexu/myalu/_0843_ ), .C1(\myexu/myalu/_1371_ ), .C2(\myexu/myalu/_0423_ ), .ZN(\myexu/myalu/_0424_ ) );
OAI21_X1 \myexu/myalu/_2689_ ( .A(\myexu/myalu/_0424_ ), .B1(\myexu/myalu/_0325_ ), .B2(\myexu/myalu/_0873_ ), .ZN(\myexu/myalu/_0425_ ) );
MUX2_X1 \myexu/myalu/_2690_ ( .A(\myexu/myalu/_0185_ ), .B(\myexu/myalu/_0425_ ), .S(\myexu/myalu/_0883_ ), .Z(\myexu/myalu/_0426_ ) );
NAND2_X1 \myexu/myalu/_2691_ ( .A1(\myexu/myalu/_0426_ ), .A2(\myexu/myalu/_0886_ ), .ZN(\myexu/myalu/_0427_ ) );
AND2_X1 \myexu/myalu/_2692_ ( .A1(\myexu/myalu/_1383_ ), .A2(\myexu/myalu/_1351_ ), .ZN(\myexu/myalu/_0429_ ) );
NAND3_X1 \myexu/myalu/_2693_ ( .A1(\myexu/myalu/_0944_ ), .A2(\myexu/myalu/_0945_ ), .A3(\myexu/myalu/_0429_ ), .ZN(\myexu/myalu/_0430_ ) );
AOI21_X1 \myexu/myalu/_2694_ ( .A(\myexu/myalu/_0872_ ), .B1(\myexu/myalu/_0557_ ), .B2(\myexu/myalu/_0753_ ), .ZN(\myexu/myalu/_0431_ ) );
AOI21_X1 \myexu/myalu/_2695_ ( .A(\myexu/myalu/_0431_ ), .B1(\myexu/myalu/_0109_ ), .B2(\myexu/myalu/_0875_ ), .ZN(\myexu/myalu/_0432_ ) );
NAND3_X1 \myexu/myalu/_2696_ ( .A1(\myexu/myalu/_0416_ ), .A2(\myexu/myalu/_0867_ ), .A3(\myexu/myalu/_0930_ ), .ZN(\myexu/myalu/_0433_ ) );
AND4_X1 \myexu/myalu/_2697_ ( .A1(\myexu/myalu/_0427_ ), .A2(\myexu/myalu/_0430_ ), .A3(\myexu/myalu/_0432_ ), .A4(\myexu/myalu/_0433_ ), .ZN(\myexu/myalu/_0434_ ) );
NAND4_X1 \myexu/myalu/_2698_ ( .A1(\myexu/myalu/_0414_ ), .A2(\myexu/myalu/_0420_ ), .A3(\myexu/myalu/_0421_ ), .A4(\myexu/myalu/_0434_ ), .ZN(\myexu/myalu/_1319_ ) );
OAI21_X1 \myexu/myalu/_2699_ ( .A(\myexu/myalu/_0220_ ), .B1(\myexu/myalu/_1287_ ), .B2(\myexu/myalu/_1292_ ), .ZN(\myexu/myalu/_0435_ ) );
MUX2_X1 \myexu/myalu/_2700_ ( .A(\myexu/myalu/_1352_ ), .B(\myexu/myalu/_1351_ ), .S(\myexu/myalu/_1360_ ), .Z(\myexu/myalu/_0436_ ) );
MUX2_X1 \myexu/myalu/_2701_ ( .A(\myexu/myalu/_0436_ ), .B(\myexu/myalu/_0399_ ), .S(\myexu/myalu/_1371_ ), .Z(\myexu/myalu/_0437_ ) );
MUX2_X1 \myexu/myalu/_2702_ ( .A(\myexu/myalu/_0437_ ), .B(\myexu/myalu/_0349_ ), .S(\myexu/myalu/_1382_ ), .Z(\myexu/myalu/_0439_ ) );
OAI21_X1 \myexu/myalu/_2703_ ( .A(\myexu/myalu/_0885_ ), .B1(\myexu/myalu/_0439_ ), .B2(\myexu/myalu/_1385_ ), .ZN(\myexu/myalu/_0440_ ) );
NOR3_X1 \myexu/myalu/_2704_ ( .A1(\myexu/myalu/_0214_ ), .A2(\myexu/myalu/_0216_ ), .A3(\myexu/myalu/_0883_ ), .ZN(\myexu/myalu/_0441_ ) );
OR2_X1 \myexu/myalu/_2705_ ( .A1(\myexu/myalu/_0440_ ), .A2(\myexu/myalu/_0441_ ), .ZN(\myexu/myalu/_0442_ ) );
AND3_X1 \myexu/myalu/_2706_ ( .A1(\myexu/myalu/_0587_ ), .A2(\myexu/myalu/_0866_ ), .A3(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_0443_ ) );
OAI21_X1 \myexu/myalu/_2707_ ( .A(\myexu/myalu/_0815_ ), .B1(\myexu/myalu/_0283_ ), .B2(\myexu/myalu/_0443_ ), .ZN(\myexu/myalu/_0444_ ) );
NAND3_X1 \myexu/myalu/_2708_ ( .A1(\myexu/myalu/_0117_ ), .A2(\myexu/myalu/_1384_ ), .A3(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_0445_ ) );
NAND4_X1 \myexu/myalu/_2709_ ( .A1(\myexu/myalu/_0587_ ), .A2(\myexu/myalu/_0866_ ), .A3(\myexu/myalu/_1352_ ), .A4(\myexu/myalu/_0929_ ), .ZN(\myexu/myalu/_0446_ ) );
NAND2_X1 \myexu/myalu/_2710_ ( .A1(\myexu/myalu/_0098_ ), .A2(\myexu/myalu/_0721_ ), .ZN(\myexu/myalu/_0447_ ) );
OAI21_X1 \myexu/myalu/_2711_ ( .A(\myexu/myalu/_0726_ ), .B1(\myexu/myalu/_1384_ ), .B2(\myexu/myalu/_1352_ ), .ZN(\myexu/myalu/_0448_ ) );
AND3_X1 \myexu/myalu/_2712_ ( .A1(\myexu/myalu/_0446_ ), .A2(\myexu/myalu/_0447_ ), .A3(\myexu/myalu/_0448_ ), .ZN(\myexu/myalu/_0450_ ) );
AND4_X1 \myexu/myalu/_2713_ ( .A1(\myexu/myalu/_0442_ ), .A2(\myexu/myalu/_0444_ ), .A3(\myexu/myalu/_0445_ ), .A4(\myexu/myalu/_0450_ ), .ZN(\myexu/myalu/_0451_ ) );
NOR2_X1 \myexu/myalu/_2714_ ( .A1(\myexu/myalu/_0412_ ), .A2(\myexu/myalu/_0429_ ), .ZN(\myexu/myalu/_0452_ ) );
XNOR2_X1 \myexu/myalu/_2715_ ( .A(\myexu/myalu/_0452_ ), .B(\myexu/myalu/_0556_ ), .ZN(\myexu/myalu/_0453_ ) );
OAI211_X2 \myexu/myalu/_2716_ ( .A(\myexu/myalu/_0435_ ), .B(\myexu/myalu/_0451_ ), .C1(\myexu/myalu/_0453_ ), .C2(\myexu/myalu/_0932_ ), .ZN(\myexu/myalu/_1320_ ) );
BUF_X1 \myexu/myalu/_2717_ ( .A(\myexu/alu_op [0] ), .Z(\myexu/myalu/_1360_ ) );
BUF_X1 \myexu/myalu/_2718_ ( .A(\src1 [0] ), .Z(\myexu/myalu/_1328_ ) );
BUF_X1 \myexu/myalu/_2719_ ( .A(\ID_EX_typ [1] ), .Z(\myexu/myalu/_0001_ ) );
BUF_X1 \myexu/myalu/_2720_ ( .A(\ID_EX_typ [0] ), .Z(\myexu/myalu/_0000_ ) );
BUF_X1 \myexu/myalu/_2721_ ( .A(\ID_EX_typ [2] ), .Z(\myexu/myalu/_0002_ ) );
BUF_X1 \myexu/myalu/_2722_ ( .A(\myexu/alu_op [4] ), .Z(\myexu/myalu/_1386_ ) );
BUF_X1 \myexu/myalu/_2723_ ( .A(\myexu/alu_op [5] ), .Z(\myexu/myalu/_1387_ ) );
BUF_X1 \myexu/myalu/_2724_ ( .A(\myexu/alu_op [3] ), .Z(\myexu/myalu/_1385_ ) );
BUF_X1 \myexu/myalu/_2725_ ( .A(\myexu/alu_op [2] ), .Z(\myexu/myalu/_1382_ ) );
BUF_X1 \myexu/myalu/_2726_ ( .A(\myexu/alu_op [1] ), .Z(\myexu/myalu/_1371_ ) );
BUF_X1 \myexu/myalu/_2727_ ( .A(\myexu/alu_op [6] ), .Z(\myexu/myalu/_1388_ ) );
BUF_X1 \myexu/myalu/_2728_ ( .A(\myexu/alu_op [7] ), .Z(\myexu/myalu/_1389_ ) );
BUF_X1 \myexu/myalu/_2729_ ( .A(\myexu/alu_op [8] ), .Z(\myexu/myalu/_1390_ ) );
BUF_X1 \myexu/myalu/_2730_ ( .A(\myexu/alu_op [9] ), .Z(\myexu/myalu/_1391_ ) );
BUF_X1 \myexu/myalu/_2731_ ( .A(\myexu/alu_op [10] ), .Z(\myexu/myalu/_1361_ ) );
BUF_X1 \myexu/myalu/_2732_ ( .A(\myexu/alu_op [11] ), .Z(\myexu/myalu/_1362_ ) );
BUF_X1 \myexu/myalu/_2733_ ( .A(\myexu/alu_op [12] ), .Z(\myexu/myalu/_1363_ ) );
BUF_X1 \myexu/myalu/_2734_ ( .A(\myexu/alu_op [13] ), .Z(\myexu/myalu/_1364_ ) );
BUF_X1 \myexu/myalu/_2735_ ( .A(\myexu/alu_op [14] ), .Z(\myexu/myalu/_1365_ ) );
BUF_X1 \myexu/myalu/_2736_ ( .A(\myexu/alu_op [15] ), .Z(\myexu/myalu/_1366_ ) );
BUF_X1 \myexu/myalu/_2737_ ( .A(\myexu/alu_op [16] ), .Z(\myexu/myalu/_1367_ ) );
BUF_X1 \myexu/myalu/_2738_ ( .A(\myexu/alu_op [17] ), .Z(\myexu/myalu/_1368_ ) );
BUF_X1 \myexu/myalu/_2739_ ( .A(\myexu/alu_op [18] ), .Z(\myexu/myalu/_1369_ ) );
BUF_X1 \myexu/myalu/_2740_ ( .A(\myexu/alu_op [19] ), .Z(\myexu/myalu/_1370_ ) );
BUF_X1 \myexu/myalu/_2741_ ( .A(\myexu/alu_op [20] ), .Z(\myexu/myalu/_1372_ ) );
BUF_X1 \myexu/myalu/_2742_ ( .A(\myexu/alu_op [21] ), .Z(\myexu/myalu/_1373_ ) );
BUF_X1 \myexu/myalu/_2743_ ( .A(\myexu/alu_op [22] ), .Z(\myexu/myalu/_1374_ ) );
BUF_X1 \myexu/myalu/_2744_ ( .A(\myexu/alu_op [23] ), .Z(\myexu/myalu/_1375_ ) );
BUF_X1 \myexu/myalu/_2745_ ( .A(\myexu/alu_op [24] ), .Z(\myexu/myalu/_1376_ ) );
BUF_X1 \myexu/myalu/_2746_ ( .A(\myexu/alu_op [25] ), .Z(\myexu/myalu/_1377_ ) );
BUF_X1 \myexu/myalu/_2747_ ( .A(\myexu/alu_op [26] ), .Z(\myexu/myalu/_1378_ ) );
BUF_X1 \myexu/myalu/_2748_ ( .A(\myexu/alu_op [27] ), .Z(\myexu/myalu/_1379_ ) );
BUF_X1 \myexu/myalu/_2749_ ( .A(\myexu/alu_op [28] ), .Z(\myexu/myalu/_1380_ ) );
BUF_X1 \myexu/myalu/_2750_ ( .A(\myexu/alu_op [29] ), .Z(\myexu/myalu/_1381_ ) );
BUF_X1 \myexu/myalu/_2751_ ( .A(\myexu/alu_op [30] ), .Z(\myexu/myalu/_1383_ ) );
BUF_X1 \myexu/myalu/_2752_ ( .A(\myexu/alu_op [31] ), .Z(\myexu/myalu/_1384_ ) );
BUF_X1 \myexu/myalu/_2753_ ( .A(\src1 [31] ), .Z(\myexu/myalu/_1352_ ) );
BUF_X1 \myexu/myalu/_2754_ ( .A(\src1 [1] ), .Z(\myexu/myalu/_1339_ ) );
BUF_X1 \myexu/myalu/_2755_ ( .A(\src1 [2] ), .Z(\myexu/myalu/_1350_ ) );
BUF_X1 \myexu/myalu/_2756_ ( .A(\src1 [3] ), .Z(\myexu/myalu/_1353_ ) );
BUF_X1 \myexu/myalu/_2757_ ( .A(\src1 [4] ), .Z(\myexu/myalu/_1354_ ) );
BUF_X1 \myexu/myalu/_2758_ ( .A(\src1 [5] ), .Z(\myexu/myalu/_1355_ ) );
BUF_X1 \myexu/myalu/_2759_ ( .A(\src1 [6] ), .Z(\myexu/myalu/_1356_ ) );
BUF_X1 \myexu/myalu/_2760_ ( .A(\src1 [7] ), .Z(\myexu/myalu/_1357_ ) );
BUF_X1 \myexu/myalu/_2761_ ( .A(\src1 [8] ), .Z(\myexu/myalu/_1358_ ) );
BUF_X1 \myexu/myalu/_2762_ ( .A(\src1 [9] ), .Z(\myexu/myalu/_1359_ ) );
BUF_X1 \myexu/myalu/_2763_ ( .A(\src1 [10] ), .Z(\myexu/myalu/_1329_ ) );
BUF_X1 \myexu/myalu/_2764_ ( .A(\src1 [11] ), .Z(\myexu/myalu/_1330_ ) );
BUF_X1 \myexu/myalu/_2765_ ( .A(\src1 [12] ), .Z(\myexu/myalu/_1331_ ) );
BUF_X1 \myexu/myalu/_2766_ ( .A(\src1 [13] ), .Z(\myexu/myalu/_1332_ ) );
BUF_X1 \myexu/myalu/_2767_ ( .A(\src1 [14] ), .Z(\myexu/myalu/_1333_ ) );
BUF_X1 \myexu/myalu/_2768_ ( .A(\src1 [15] ), .Z(\myexu/myalu/_1334_ ) );
BUF_X1 \myexu/myalu/_2769_ ( .A(\src1 [16] ), .Z(\myexu/myalu/_1335_ ) );
BUF_X1 \myexu/myalu/_2770_ ( .A(\src1 [17] ), .Z(\myexu/myalu/_1336_ ) );
BUF_X1 \myexu/myalu/_2771_ ( .A(\src1 [18] ), .Z(\myexu/myalu/_1337_ ) );
BUF_X1 \myexu/myalu/_2772_ ( .A(\src1 [19] ), .Z(\myexu/myalu/_1338_ ) );
BUF_X1 \myexu/myalu/_2773_ ( .A(\src1 [20] ), .Z(\myexu/myalu/_1340_ ) );
BUF_X1 \myexu/myalu/_2774_ ( .A(\src1 [21] ), .Z(\myexu/myalu/_1341_ ) );
BUF_X1 \myexu/myalu/_2775_ ( .A(\src1 [22] ), .Z(\myexu/myalu/_1342_ ) );
BUF_X1 \myexu/myalu/_2776_ ( .A(\src1 [23] ), .Z(\myexu/myalu/_1343_ ) );
BUF_X1 \myexu/myalu/_2777_ ( .A(\src1 [24] ), .Z(\myexu/myalu/_1344_ ) );
BUF_X1 \myexu/myalu/_2778_ ( .A(\src1 [25] ), .Z(\myexu/myalu/_1345_ ) );
BUF_X1 \myexu/myalu/_2779_ ( .A(\src1 [26] ), .Z(\myexu/myalu/_1346_ ) );
BUF_X1 \myexu/myalu/_2780_ ( .A(\src1 [27] ), .Z(\myexu/myalu/_1347_ ) );
BUF_X1 \myexu/myalu/_2781_ ( .A(\src1 [28] ), .Z(\myexu/myalu/_1348_ ) );
BUF_X1 \myexu/myalu/_2782_ ( .A(\src1 [29] ), .Z(\myexu/myalu/_1349_ ) );
BUF_X1 \myexu/myalu/_2783_ ( .A(\src1 [30] ), .Z(\myexu/myalu/_1351_ ) );
BUF_X1 \myexu/myalu/_2784_ ( .A(\myexu/myalu/_1296_ ), .Z(\myexu/alu_out [0] ) );
BUF_X1 \myexu/myalu/_2785_ ( .A(\myexu/myalu/_1307_ ), .Z(\myexu/alu_out [1] ) );
BUF_X1 \myexu/myalu/_2786_ ( .A(\myexu/myalu/_1318_ ), .Z(\myexu/alu_out [2] ) );
BUF_X1 \myexu/myalu/_2787_ ( .A(\myexu/myalu/_1321_ ), .Z(\myexu/alu_out [3] ) );
BUF_X1 \myexu/myalu/_2788_ ( .A(\myexu/myalu/_1322_ ), .Z(\myexu/alu_out [4] ) );
BUF_X1 \myexu/myalu/_2789_ ( .A(\myexu/myalu/_1323_ ), .Z(\myexu/alu_out [5] ) );
BUF_X1 \myexu/myalu/_2790_ ( .A(\myexu/myalu/_1324_ ), .Z(\myexu/alu_out [6] ) );
BUF_X1 \myexu/myalu/_2791_ ( .A(\myexu/myalu/_1325_ ), .Z(\myexu/alu_out [7] ) );
BUF_X1 \myexu/myalu/_2792_ ( .A(\myexu/myalu/_1326_ ), .Z(\myexu/alu_out [8] ) );
BUF_X1 \myexu/myalu/_2793_ ( .A(\myexu/myalu/_1327_ ), .Z(\myexu/alu_out [9] ) );
BUF_X1 \myexu/myalu/_2794_ ( .A(\myexu/myalu/_1297_ ), .Z(\myexu/alu_out [10] ) );
BUF_X1 \myexu/myalu/_2795_ ( .A(\myexu/myalu/_1298_ ), .Z(\myexu/alu_out [11] ) );
BUF_X1 \myexu/myalu/_2796_ ( .A(\myexu/myalu/_1299_ ), .Z(\myexu/alu_out [12] ) );
BUF_X1 \myexu/myalu/_2797_ ( .A(\myexu/myalu/_1300_ ), .Z(\myexu/alu_out [13] ) );
BUF_X1 \myexu/myalu/_2798_ ( .A(\myexu/myalu/_1301_ ), .Z(\myexu/alu_out [14] ) );
BUF_X1 \myexu/myalu/_2799_ ( .A(\myexu/myalu/_1302_ ), .Z(\myexu/alu_out [15] ) );
BUF_X1 \myexu/myalu/_2800_ ( .A(\myexu/myalu/_1303_ ), .Z(\myexu/alu_out [16] ) );
BUF_X1 \myexu/myalu/_2801_ ( .A(\myexu/myalu/_1304_ ), .Z(\myexu/alu_out [17] ) );
BUF_X1 \myexu/myalu/_2802_ ( .A(\myexu/myalu/_1305_ ), .Z(\myexu/alu_out [18] ) );
BUF_X1 \myexu/myalu/_2803_ ( .A(\myexu/myalu/_1306_ ), .Z(\myexu/alu_out [19] ) );
BUF_X1 \myexu/myalu/_2804_ ( .A(\myexu/myalu/_1308_ ), .Z(\myexu/alu_out [20] ) );
BUF_X1 \myexu/myalu/_2805_ ( .A(\myexu/myalu/_1309_ ), .Z(\myexu/alu_out [21] ) );
BUF_X1 \myexu/myalu/_2806_ ( .A(\myexu/myalu/_1310_ ), .Z(\myexu/alu_out [22] ) );
BUF_X1 \myexu/myalu/_2807_ ( .A(\myexu/myalu/_1311_ ), .Z(\myexu/alu_out [23] ) );
BUF_X1 \myexu/myalu/_2808_ ( .A(\myexu/myalu/_1312_ ), .Z(\myexu/alu_out [24] ) );
BUF_X1 \myexu/myalu/_2809_ ( .A(\myexu/myalu/_1313_ ), .Z(\myexu/alu_out [25] ) );
BUF_X1 \myexu/myalu/_2810_ ( .A(\myexu/myalu/_1314_ ), .Z(\myexu/alu_out [26] ) );
BUF_X1 \myexu/myalu/_2811_ ( .A(\myexu/myalu/_1315_ ), .Z(\myexu/alu_out [27] ) );
BUF_X1 \myexu/myalu/_2812_ ( .A(\myexu/myalu/_1316_ ), .Z(\myexu/alu_out [28] ) );
BUF_X1 \myexu/myalu/_2813_ ( .A(\myexu/myalu/_1317_ ), .Z(\myexu/alu_out [29] ) );
BUF_X1 \myexu/myalu/_2814_ ( .A(\myexu/myalu/_1319_ ), .Z(\myexu/alu_out [30] ) );
BUF_X1 \myexu/myalu/_2815_ ( .A(\myexu/myalu/_1320_ ), .Z(\myexu/alu_out [31] ) );
OR4_X1 \myfc/_385_ ( .A1(\myfc/_014_ ), .A2(\myfc/_015_ ), .A3(\myfc/_016_ ), .A4(\myfc/_017_ ), .ZN(\myfc/_138_ ) );
OR2_X1 \myfc/_386_ ( .A1(\myfc/_138_ ), .A2(\myfc/_018_ ), .ZN(\myfc/_139_ ) );
XNOR2_X1 \myfc/_387_ ( .A(\myfc/_031_ ), .B(\myfc/_014_ ), .ZN(\myfc/_140_ ) );
XNOR2_X1 \myfc/_388_ ( .A(\myfc/_033_ ), .B(\myfc/_016_ ), .ZN(\myfc/_141_ ) );
XNOR2_X1 \myfc/_389_ ( .A(\myfc/_034_ ), .B(\myfc/_017_ ), .ZN(\myfc/_142_ ) );
XNOR2_X1 \myfc/_390_ ( .A(\myfc/_032_ ), .B(\myfc/_015_ ), .ZN(\myfc/_143_ ) );
AND4_X1 \myfc/_391_ ( .A1(\myfc/_140_ ), .A2(\myfc/_141_ ), .A3(\myfc/_142_ ), .A4(\myfc/_143_ ), .ZN(\myfc/_144_ ) );
XNOR2_X1 \myfc/_392_ ( .A(\myfc/_035_ ), .B(\myfc/_018_ ), .ZN(\myfc/_145_ ) );
NAND4_X1 \myfc/_393_ ( .A1(\myfc/_139_ ), .A2(\myfc/_144_ ), .A3(\myfc/_001_ ), .A4(\myfc/_145_ ), .ZN(\myfc/_146_ ) );
NOR2_X1 \myfc/_394_ ( .A1(\myfc/_146_ ), .A2(\myfc/_137_ ), .ZN(\myfc/_147_ ) );
BUF_X4 \myfc/_395_ ( .A(\myfc/_147_ ), .Z(\myfc/_148_ ) );
MUX2_X1 \myfc/_396_ ( .A(\myfc/_193_ ), .B(\myfc/_041_ ), .S(\myfc/_148_ ), .Z(\myfc/_289_ ) );
MUX2_X1 \myfc/_397_ ( .A(\myfc/_204_ ), .B(\myfc/_052_ ), .S(\myfc/_148_ ), .Z(\myfc/_300_ ) );
MUX2_X1 \myfc/_398_ ( .A(\myfc/_215_ ), .B(\myfc/_063_ ), .S(\myfc/_148_ ), .Z(\myfc/_311_ ) );
MUX2_X1 \myfc/_399_ ( .A(\myfc/_218_ ), .B(\myfc/_066_ ), .S(\myfc/_148_ ), .Z(\myfc/_314_ ) );
MUX2_X1 \myfc/_400_ ( .A(\myfc/_219_ ), .B(\myfc/_067_ ), .S(\myfc/_148_ ), .Z(\myfc/_315_ ) );
MUX2_X1 \myfc/_401_ ( .A(\myfc/_220_ ), .B(\myfc/_068_ ), .S(\myfc/_148_ ), .Z(\myfc/_316_ ) );
MUX2_X1 \myfc/_402_ ( .A(\myfc/_221_ ), .B(\myfc/_069_ ), .S(\myfc/_148_ ), .Z(\myfc/_317_ ) );
MUX2_X1 \myfc/_403_ ( .A(\myfc/_222_ ), .B(\myfc/_070_ ), .S(\myfc/_148_ ), .Z(\myfc/_318_ ) );
MUX2_X1 \myfc/_404_ ( .A(\myfc/_223_ ), .B(\myfc/_071_ ), .S(\myfc/_148_ ), .Z(\myfc/_319_ ) );
MUX2_X1 \myfc/_405_ ( .A(\myfc/_224_ ), .B(\myfc/_072_ ), .S(\myfc/_148_ ), .Z(\myfc/_320_ ) );
BUF_X4 \myfc/_406_ ( .A(\myfc/_147_ ), .Z(\myfc/_149_ ) );
MUX2_X1 \myfc/_407_ ( .A(\myfc/_194_ ), .B(\myfc/_042_ ), .S(\myfc/_149_ ), .Z(\myfc/_290_ ) );
MUX2_X1 \myfc/_408_ ( .A(\myfc/_195_ ), .B(\myfc/_043_ ), .S(\myfc/_149_ ), .Z(\myfc/_291_ ) );
MUX2_X1 \myfc/_409_ ( .A(\myfc/_196_ ), .B(\myfc/_044_ ), .S(\myfc/_149_ ), .Z(\myfc/_292_ ) );
MUX2_X1 \myfc/_410_ ( .A(\myfc/_197_ ), .B(\myfc/_045_ ), .S(\myfc/_149_ ), .Z(\myfc/_293_ ) );
MUX2_X1 \myfc/_411_ ( .A(\myfc/_198_ ), .B(\myfc/_046_ ), .S(\myfc/_149_ ), .Z(\myfc/_294_ ) );
MUX2_X1 \myfc/_412_ ( .A(\myfc/_199_ ), .B(\myfc/_047_ ), .S(\myfc/_149_ ), .Z(\myfc/_295_ ) );
MUX2_X1 \myfc/_413_ ( .A(\myfc/_200_ ), .B(\myfc/_048_ ), .S(\myfc/_149_ ), .Z(\myfc/_296_ ) );
MUX2_X1 \myfc/_414_ ( .A(\myfc/_201_ ), .B(\myfc/_049_ ), .S(\myfc/_149_ ), .Z(\myfc/_297_ ) );
MUX2_X1 \myfc/_415_ ( .A(\myfc/_202_ ), .B(\myfc/_050_ ), .S(\myfc/_149_ ), .Z(\myfc/_298_ ) );
MUX2_X1 \myfc/_416_ ( .A(\myfc/_203_ ), .B(\myfc/_051_ ), .S(\myfc/_149_ ), .Z(\myfc/_299_ ) );
BUF_X4 \myfc/_417_ ( .A(\myfc/_147_ ), .Z(\myfc/_150_ ) );
MUX2_X1 \myfc/_418_ ( .A(\myfc/_205_ ), .B(\myfc/_053_ ), .S(\myfc/_150_ ), .Z(\myfc/_301_ ) );
MUX2_X1 \myfc/_419_ ( .A(\myfc/_206_ ), .B(\myfc/_054_ ), .S(\myfc/_150_ ), .Z(\myfc/_302_ ) );
MUX2_X1 \myfc/_420_ ( .A(\myfc/_207_ ), .B(\myfc/_055_ ), .S(\myfc/_150_ ), .Z(\myfc/_303_ ) );
MUX2_X1 \myfc/_421_ ( .A(\myfc/_208_ ), .B(\myfc/_056_ ), .S(\myfc/_150_ ), .Z(\myfc/_304_ ) );
MUX2_X1 \myfc/_422_ ( .A(\myfc/_209_ ), .B(\myfc/_057_ ), .S(\myfc/_150_ ), .Z(\myfc/_305_ ) );
MUX2_X1 \myfc/_423_ ( .A(\myfc/_210_ ), .B(\myfc/_058_ ), .S(\myfc/_150_ ), .Z(\myfc/_306_ ) );
MUX2_X1 \myfc/_424_ ( .A(\myfc/_211_ ), .B(\myfc/_059_ ), .S(\myfc/_150_ ), .Z(\myfc/_307_ ) );
MUX2_X1 \myfc/_425_ ( .A(\myfc/_212_ ), .B(\myfc/_060_ ), .S(\myfc/_150_ ), .Z(\myfc/_308_ ) );
MUX2_X1 \myfc/_426_ ( .A(\myfc/_213_ ), .B(\myfc/_061_ ), .S(\myfc/_150_ ), .Z(\myfc/_309_ ) );
MUX2_X1 \myfc/_427_ ( .A(\myfc/_214_ ), .B(\myfc/_062_ ), .S(\myfc/_150_ ), .Z(\myfc/_310_ ) );
MUX2_X1 \myfc/_428_ ( .A(\myfc/_216_ ), .B(\myfc/_064_ ), .S(\myfc/_147_ ), .Z(\myfc/_312_ ) );
MUX2_X1 \myfc/_429_ ( .A(\myfc/_217_ ), .B(\myfc/_065_ ), .S(\myfc/_147_ ), .Z(\myfc/_313_ ) );
XNOR2_X1 \myfc/_430_ ( .A(\myfc/_014_ ), .B(\myfc/_036_ ), .ZN(\myfc/_151_ ) );
XNOR2_X1 \myfc/_431_ ( .A(\myfc/_016_ ), .B(\myfc/_038_ ), .ZN(\myfc/_152_ ) );
XNOR2_X1 \myfc/_432_ ( .A(\myfc/_017_ ), .B(\myfc/_039_ ), .ZN(\myfc/_153_ ) );
XNOR2_X1 \myfc/_433_ ( .A(\myfc/_015_ ), .B(\myfc/_037_ ), .ZN(\myfc/_154_ ) );
AND4_X1 \myfc/_434_ ( .A1(\myfc/_151_ ), .A2(\myfc/_152_ ), .A3(\myfc/_153_ ), .A4(\myfc/_154_ ), .ZN(\myfc/_155_ ) );
XNOR2_X1 \myfc/_435_ ( .A(\myfc/_018_ ), .B(\myfc/_040_ ), .ZN(\myfc/_156_ ) );
NAND4_X1 \myfc/_436_ ( .A1(\myfc/_139_ ), .A2(\myfc/_155_ ), .A3(\myfc/_001_ ), .A4(\myfc/_156_ ), .ZN(\myfc/_157_ ) );
NOR2_X1 \myfc/_437_ ( .A1(\myfc/_157_ ), .A2(\myfc/_137_ ), .ZN(\myfc/_158_ ) );
BUF_X4 \myfc/_438_ ( .A(\myfc/_158_ ), .Z(\myfc/_159_ ) );
MUX2_X1 \myfc/_439_ ( .A(\myfc/_225_ ), .B(\myfc/_073_ ), .S(\myfc/_159_ ), .Z(\myfc/_321_ ) );
MUX2_X1 \myfc/_440_ ( .A(\myfc/_236_ ), .B(\myfc/_084_ ), .S(\myfc/_159_ ), .Z(\myfc/_332_ ) );
MUX2_X1 \myfc/_441_ ( .A(\myfc/_247_ ), .B(\myfc/_095_ ), .S(\myfc/_159_ ), .Z(\myfc/_343_ ) );
MUX2_X1 \myfc/_442_ ( .A(\myfc/_250_ ), .B(\myfc/_098_ ), .S(\myfc/_159_ ), .Z(\myfc/_346_ ) );
MUX2_X1 \myfc/_443_ ( .A(\myfc/_251_ ), .B(\myfc/_099_ ), .S(\myfc/_159_ ), .Z(\myfc/_347_ ) );
MUX2_X1 \myfc/_444_ ( .A(\myfc/_252_ ), .B(\myfc/_100_ ), .S(\myfc/_159_ ), .Z(\myfc/_348_ ) );
MUX2_X1 \myfc/_445_ ( .A(\myfc/_253_ ), .B(\myfc/_101_ ), .S(\myfc/_159_ ), .Z(\myfc/_349_ ) );
MUX2_X1 \myfc/_446_ ( .A(\myfc/_254_ ), .B(\myfc/_102_ ), .S(\myfc/_159_ ), .Z(\myfc/_350_ ) );
MUX2_X1 \myfc/_447_ ( .A(\myfc/_255_ ), .B(\myfc/_103_ ), .S(\myfc/_159_ ), .Z(\myfc/_351_ ) );
MUX2_X1 \myfc/_448_ ( .A(\myfc/_256_ ), .B(\myfc/_104_ ), .S(\myfc/_159_ ), .Z(\myfc/_352_ ) );
BUF_X4 \myfc/_449_ ( .A(\myfc/_158_ ), .Z(\myfc/_160_ ) );
MUX2_X1 \myfc/_450_ ( .A(\myfc/_226_ ), .B(\myfc/_074_ ), .S(\myfc/_160_ ), .Z(\myfc/_322_ ) );
MUX2_X1 \myfc/_451_ ( .A(\myfc/_227_ ), .B(\myfc/_075_ ), .S(\myfc/_160_ ), .Z(\myfc/_323_ ) );
MUX2_X1 \myfc/_452_ ( .A(\myfc/_228_ ), .B(\myfc/_076_ ), .S(\myfc/_160_ ), .Z(\myfc/_324_ ) );
MUX2_X1 \myfc/_453_ ( .A(\myfc/_229_ ), .B(\myfc/_077_ ), .S(\myfc/_160_ ), .Z(\myfc/_325_ ) );
MUX2_X1 \myfc/_454_ ( .A(\myfc/_230_ ), .B(\myfc/_078_ ), .S(\myfc/_160_ ), .Z(\myfc/_326_ ) );
MUX2_X1 \myfc/_455_ ( .A(\myfc/_231_ ), .B(\myfc/_079_ ), .S(\myfc/_160_ ), .Z(\myfc/_327_ ) );
MUX2_X1 \myfc/_456_ ( .A(\myfc/_232_ ), .B(\myfc/_080_ ), .S(\myfc/_160_ ), .Z(\myfc/_328_ ) );
MUX2_X1 \myfc/_457_ ( .A(\myfc/_233_ ), .B(\myfc/_081_ ), .S(\myfc/_160_ ), .Z(\myfc/_329_ ) );
MUX2_X1 \myfc/_458_ ( .A(\myfc/_234_ ), .B(\myfc/_082_ ), .S(\myfc/_160_ ), .Z(\myfc/_330_ ) );
MUX2_X1 \myfc/_459_ ( .A(\myfc/_235_ ), .B(\myfc/_083_ ), .S(\myfc/_160_ ), .Z(\myfc/_331_ ) );
BUF_X4 \myfc/_460_ ( .A(\myfc/_158_ ), .Z(\myfc/_161_ ) );
MUX2_X1 \myfc/_461_ ( .A(\myfc/_237_ ), .B(\myfc/_085_ ), .S(\myfc/_161_ ), .Z(\myfc/_333_ ) );
MUX2_X1 \myfc/_462_ ( .A(\myfc/_238_ ), .B(\myfc/_086_ ), .S(\myfc/_161_ ), .Z(\myfc/_334_ ) );
MUX2_X1 \myfc/_463_ ( .A(\myfc/_239_ ), .B(\myfc/_087_ ), .S(\myfc/_161_ ), .Z(\myfc/_335_ ) );
MUX2_X1 \myfc/_464_ ( .A(\myfc/_240_ ), .B(\myfc/_088_ ), .S(\myfc/_161_ ), .Z(\myfc/_336_ ) );
MUX2_X1 \myfc/_465_ ( .A(\myfc/_241_ ), .B(\myfc/_089_ ), .S(\myfc/_161_ ), .Z(\myfc/_337_ ) );
MUX2_X1 \myfc/_466_ ( .A(\myfc/_242_ ), .B(\myfc/_090_ ), .S(\myfc/_161_ ), .Z(\myfc/_338_ ) );
MUX2_X1 \myfc/_467_ ( .A(\myfc/_243_ ), .B(\myfc/_091_ ), .S(\myfc/_161_ ), .Z(\myfc/_339_ ) );
MUX2_X1 \myfc/_468_ ( .A(\myfc/_244_ ), .B(\myfc/_092_ ), .S(\myfc/_161_ ), .Z(\myfc/_340_ ) );
MUX2_X1 \myfc/_469_ ( .A(\myfc/_245_ ), .B(\myfc/_093_ ), .S(\myfc/_161_ ), .Z(\myfc/_341_ ) );
MUX2_X1 \myfc/_470_ ( .A(\myfc/_246_ ), .B(\myfc/_094_ ), .S(\myfc/_161_ ), .Z(\myfc/_342_ ) );
MUX2_X1 \myfc/_471_ ( .A(\myfc/_248_ ), .B(\myfc/_096_ ), .S(\myfc/_158_ ), .Z(\myfc/_344_ ) );
MUX2_X1 \myfc/_472_ ( .A(\myfc/_249_ ), .B(\myfc/_097_ ), .S(\myfc/_158_ ), .Z(\myfc/_345_ ) );
XOR2_X2 \myfc/_473_ ( .A(\myfc/_029_ ), .B(\myfc/_012_ ), .Z(\myfc/_162_ ) );
INV_X1 \myfc/_474_ ( .A(\myfc/_028_ ), .ZN(\myfc/_163_ ) );
AND2_X1 \myfc/_475_ ( .A1(\myfc/_163_ ), .A2(\myfc/_011_ ), .ZN(\myfc/_164_ ) );
INV_X1 \myfc/_476_ ( .A(\myfc/_030_ ), .ZN(\myfc/_165_ ) );
NOR2_X1 \myfc/_477_ ( .A1(\myfc/_165_ ), .A2(\myfc/_013_ ), .ZN(\myfc/_166_ ) );
OR3_X4 \myfc/_478_ ( .A1(\myfc/_162_ ), .A2(\myfc/_164_ ), .A3(\myfc/_166_ ), .ZN(\myfc/_167_ ) );
INV_X1 \myfc/_479_ ( .A(\myfc/_004_ ), .ZN(\myfc/_168_ ) );
AOI221_X2 \myfc/_480_ ( .A(\myfc/_167_ ), .B1(\myfc/_165_ ), .B2(\myfc/_013_ ), .C1(\myfc/_021_ ), .C2(\myfc/_168_ ), .ZN(\myfc/_169_ ) );
INV_X1 \myfc/_481_ ( .A(\myfc/_002_ ), .ZN(\myfc/_170_ ) );
OR2_X1 \myfc/_482_ ( .A1(\myfc/_170_ ), .A2(\myfc/_019_ ), .ZN(\myfc/_171_ ) );
INV_X1 \myfc/_483_ ( .A(\myfc/_005_ ), .ZN(\myfc/_172_ ) );
AOI22_X1 \myfc/_484_ ( .A1(\myfc/_019_ ), .A2(\myfc/_170_ ), .B1(\myfc/_172_ ), .B2(\myfc/_022_ ), .ZN(\myfc/_173_ ) );
INV_X1 \myfc/_485_ ( .A(\myfc/_026_ ), .ZN(\myfc/_174_ ) );
NOR2_X1 \myfc/_486_ ( .A1(\myfc/_174_ ), .A2(\myfc/_009_ ), .ZN(\myfc/_175_ ) );
INV_X1 \myfc/_487_ ( .A(\myfc/_024_ ), .ZN(\myfc/_176_ ) );
OAI22_X1 \myfc/_488_ ( .A1(\myfc/_022_ ), .A2(\myfc/_172_ ), .B1(\myfc/_176_ ), .B2(\myfc/_007_ ), .ZN(\myfc/_177_ ) );
AOI211_X4 \myfc/_489_ ( .A(\myfc/_175_ ), .B(\myfc/_177_ ), .C1(\myfc/_176_ ), .C2(\myfc/_007_ ), .ZN(\myfc/_178_ ) );
NAND4_X2 \myfc/_490_ ( .A1(\myfc/_169_ ), .A2(\myfc/_171_ ), .A3(\myfc/_173_ ), .A4(\myfc/_178_ ), .ZN(\myfc/_179_ ) );
NOR2_X1 \myfc/_491_ ( .A1(\myfc/_163_ ), .A2(\myfc/_011_ ), .ZN(\myfc/_180_ ) );
XOR2_X1 \myfc/_492_ ( .A(\myfc/_027_ ), .B(\myfc/_010_ ), .Z(\myfc/_181_ ) );
AOI211_X4 \myfc/_493_ ( .A(\myfc/_180_ ), .B(\myfc/_181_ ), .C1(\myfc/_174_ ), .C2(\myfc/_009_ ), .ZN(\myfc/_182_ ) );
XNOR2_X1 \myfc/_494_ ( .A(\myfc/_020_ ), .B(\myfc/_003_ ), .ZN(\myfc/_183_ ) );
OR2_X1 \myfc/_495_ ( .A1(\myfc/_168_ ), .A2(\myfc/_021_ ), .ZN(\myfc/_184_ ) );
AND3_X1 \myfc/_496_ ( .A1(\myfc/_183_ ), .A2(\myfc/_000_ ), .A3(\myfc/_184_ ), .ZN(\myfc/_185_ ) );
XNOR2_X1 \myfc/_497_ ( .A(\myfc/_025_ ), .B(\myfc/_008_ ), .ZN(\myfc/_186_ ) );
XNOR2_X1 \myfc/_498_ ( .A(\myfc/_023_ ), .B(\myfc/_006_ ), .ZN(\myfc/_187_ ) );
NAND4_X1 \myfc/_499_ ( .A1(\myfc/_182_ ), .A2(\myfc/_185_ ), .A3(\myfc/_186_ ), .A4(\myfc/_187_ ), .ZN(\myfc/_188_ ) );
NOR2_X4 \myfc/_500_ ( .A1(\myfc/_179_ ), .A2(\myfc/_188_ ), .ZN(\myfc/_189_ ) );
BUF_X4 \myfc/_501_ ( .A(\myfc/_189_ ), .Z(\myfc/_190_ ) );
MUX2_X1 \myfc/_502_ ( .A(\myfc/_257_ ), .B(\myfc/_105_ ), .S(\myfc/_190_ ), .Z(\myfc/_353_ ) );
MUX2_X1 \myfc/_503_ ( .A(\myfc/_268_ ), .B(\myfc/_116_ ), .S(\myfc/_190_ ), .Z(\myfc/_364_ ) );
MUX2_X1 \myfc/_504_ ( .A(\myfc/_279_ ), .B(\myfc/_127_ ), .S(\myfc/_190_ ), .Z(\myfc/_375_ ) );
MUX2_X1 \myfc/_505_ ( .A(\myfc/_282_ ), .B(\myfc/_130_ ), .S(\myfc/_190_ ), .Z(\myfc/_378_ ) );
MUX2_X1 \myfc/_506_ ( .A(\myfc/_283_ ), .B(\myfc/_131_ ), .S(\myfc/_190_ ), .Z(\myfc/_379_ ) );
MUX2_X1 \myfc/_507_ ( .A(\myfc/_284_ ), .B(\myfc/_132_ ), .S(\myfc/_190_ ), .Z(\myfc/_380_ ) );
MUX2_X1 \myfc/_508_ ( .A(\myfc/_285_ ), .B(\myfc/_133_ ), .S(\myfc/_190_ ), .Z(\myfc/_381_ ) );
MUX2_X1 \myfc/_509_ ( .A(\myfc/_286_ ), .B(\myfc/_134_ ), .S(\myfc/_190_ ), .Z(\myfc/_382_ ) );
MUX2_X1 \myfc/_510_ ( .A(\myfc/_287_ ), .B(\myfc/_135_ ), .S(\myfc/_190_ ), .Z(\myfc/_383_ ) );
MUX2_X1 \myfc/_511_ ( .A(\myfc/_288_ ), .B(\myfc/_136_ ), .S(\myfc/_190_ ), .Z(\myfc/_384_ ) );
BUF_X8 \myfc/_512_ ( .A(\myfc/_189_ ), .Z(\myfc/_191_ ) );
MUX2_X1 \myfc/_513_ ( .A(\myfc/_258_ ), .B(\myfc/_106_ ), .S(\myfc/_191_ ), .Z(\myfc/_354_ ) );
MUX2_X1 \myfc/_514_ ( .A(\myfc/_259_ ), .B(\myfc/_107_ ), .S(\myfc/_191_ ), .Z(\myfc/_355_ ) );
MUX2_X1 \myfc/_515_ ( .A(\myfc/_260_ ), .B(\myfc/_108_ ), .S(\myfc/_191_ ), .Z(\myfc/_356_ ) );
MUX2_X1 \myfc/_516_ ( .A(\myfc/_261_ ), .B(\myfc/_109_ ), .S(\myfc/_191_ ), .Z(\myfc/_357_ ) );
MUX2_X1 \myfc/_517_ ( .A(\myfc/_262_ ), .B(\myfc/_110_ ), .S(\myfc/_191_ ), .Z(\myfc/_358_ ) );
MUX2_X1 \myfc/_518_ ( .A(\myfc/_263_ ), .B(\myfc/_111_ ), .S(\myfc/_191_ ), .Z(\myfc/_359_ ) );
MUX2_X1 \myfc/_519_ ( .A(\myfc/_264_ ), .B(\myfc/_112_ ), .S(\myfc/_191_ ), .Z(\myfc/_360_ ) );
MUX2_X1 \myfc/_520_ ( .A(\myfc/_265_ ), .B(\myfc/_113_ ), .S(\myfc/_191_ ), .Z(\myfc/_361_ ) );
MUX2_X1 \myfc/_521_ ( .A(\myfc/_266_ ), .B(\myfc/_114_ ), .S(\myfc/_191_ ), .Z(\myfc/_362_ ) );
MUX2_X1 \myfc/_522_ ( .A(\myfc/_267_ ), .B(\myfc/_115_ ), .S(\myfc/_191_ ), .Z(\myfc/_363_ ) );
BUF_X4 \myfc/_523_ ( .A(\myfc/_189_ ), .Z(\myfc/_192_ ) );
MUX2_X1 \myfc/_524_ ( .A(\myfc/_269_ ), .B(\myfc/_117_ ), .S(\myfc/_192_ ), .Z(\myfc/_365_ ) );
MUX2_X1 \myfc/_525_ ( .A(\myfc/_270_ ), .B(\myfc/_118_ ), .S(\myfc/_192_ ), .Z(\myfc/_366_ ) );
MUX2_X1 \myfc/_526_ ( .A(\myfc/_271_ ), .B(\myfc/_119_ ), .S(\myfc/_192_ ), .Z(\myfc/_367_ ) );
MUX2_X1 \myfc/_527_ ( .A(\myfc/_272_ ), .B(\myfc/_120_ ), .S(\myfc/_192_ ), .Z(\myfc/_368_ ) );
MUX2_X1 \myfc/_528_ ( .A(\myfc/_273_ ), .B(\myfc/_121_ ), .S(\myfc/_192_ ), .Z(\myfc/_369_ ) );
MUX2_X1 \myfc/_529_ ( .A(\myfc/_274_ ), .B(\myfc/_122_ ), .S(\myfc/_192_ ), .Z(\myfc/_370_ ) );
MUX2_X1 \myfc/_530_ ( .A(\myfc/_275_ ), .B(\myfc/_123_ ), .S(\myfc/_192_ ), .Z(\myfc/_371_ ) );
MUX2_X1 \myfc/_531_ ( .A(\myfc/_276_ ), .B(\myfc/_124_ ), .S(\myfc/_192_ ), .Z(\myfc/_372_ ) );
MUX2_X1 \myfc/_532_ ( .A(\myfc/_277_ ), .B(\myfc/_125_ ), .S(\myfc/_192_ ), .Z(\myfc/_373_ ) );
MUX2_X1 \myfc/_533_ ( .A(\myfc/_278_ ), .B(\myfc/_126_ ), .S(\myfc/_192_ ), .Z(\myfc/_374_ ) );
MUX2_X1 \myfc/_534_ ( .A(\myfc/_280_ ), .B(\myfc/_128_ ), .S(\myfc/_189_ ), .Z(\myfc/_376_ ) );
MUX2_X1 \myfc/_535_ ( .A(\myfc/_281_ ), .B(\myfc/_129_ ), .S(\myfc/_189_ ), .Z(\myfc/_377_ ) );
BUF_X1 \myfc/_536_ ( .A(EX_LS_RegWrite ), .Z(\myfc/_001_ ) );
BUF_X1 \myfc/_537_ ( .A(\ID_EX_rs1 [0] ), .Z(\myfc/_031_ ) );
BUF_X1 \myfc/_538_ ( .A(\EX_LS_dest_reg [0] ), .Z(\myfc/_014_ ) );
BUF_X1 \myfc/_539_ ( .A(\ID_EX_rs1 [1] ), .Z(\myfc/_032_ ) );
BUF_X1 \myfc/_540_ ( .A(\EX_LS_dest_reg [1] ), .Z(\myfc/_015_ ) );
BUF_X1 \myfc/_541_ ( .A(\ID_EX_rs1 [2] ), .Z(\myfc/_033_ ) );
BUF_X1 \myfc/_542_ ( .A(\EX_LS_dest_reg [2] ), .Z(\myfc/_016_ ) );
BUF_X1 \myfc/_543_ ( .A(\ID_EX_rs1 [3] ), .Z(\myfc/_034_ ) );
BUF_X1 \myfc/_544_ ( .A(\EX_LS_dest_reg [3] ), .Z(\myfc/_017_ ) );
BUF_X1 \myfc/_545_ ( .A(\ID_EX_rs1 [4] ), .Z(\myfc/_035_ ) );
BUF_X1 \myfc/_546_ ( .A(\EX_LS_dest_reg [4] ), .Z(\myfc/_018_ ) );
BUF_X1 \myfc/_547_ ( .A(fc_disenable ), .Z(\myfc/_137_ ) );
BUF_X1 \myfc/_548_ ( .A(\EX_LS_result_reg [0] ), .Z(\myfc/_041_ ) );
BUF_X1 \myfc/_549_ ( .A(\src1_raw [0] ), .Z(\myfc/_193_ ) );
BUF_X1 \myfc/_550_ ( .A(\myfc/_289_ ), .Z(\src1 [0] ) );
BUF_X1 \myfc/_551_ ( .A(\EX_LS_result_reg [1] ), .Z(\myfc/_052_ ) );
BUF_X1 \myfc/_552_ ( .A(\src1_raw [1] ), .Z(\myfc/_204_ ) );
BUF_X1 \myfc/_553_ ( .A(\myfc/_300_ ), .Z(\src1 [1] ) );
BUF_X1 \myfc/_554_ ( .A(\EX_LS_result_reg [2] ), .Z(\myfc/_063_ ) );
BUF_X1 \myfc/_555_ ( .A(\src1_raw [2] ), .Z(\myfc/_215_ ) );
BUF_X1 \myfc/_556_ ( .A(\myfc/_311_ ), .Z(\src1 [2] ) );
BUF_X1 \myfc/_557_ ( .A(\EX_LS_result_reg [3] ), .Z(\myfc/_066_ ) );
BUF_X1 \myfc/_558_ ( .A(\src1_raw [3] ), .Z(\myfc/_218_ ) );
BUF_X1 \myfc/_559_ ( .A(\myfc/_314_ ), .Z(\src1 [3] ) );
BUF_X1 \myfc/_560_ ( .A(\EX_LS_result_reg [4] ), .Z(\myfc/_067_ ) );
BUF_X1 \myfc/_561_ ( .A(\src1_raw [4] ), .Z(\myfc/_219_ ) );
BUF_X1 \myfc/_562_ ( .A(\myfc/_315_ ), .Z(\src1 [4] ) );
BUF_X1 \myfc/_563_ ( .A(\EX_LS_result_reg [5] ), .Z(\myfc/_068_ ) );
BUF_X1 \myfc/_564_ ( .A(\src1_raw [5] ), .Z(\myfc/_220_ ) );
BUF_X1 \myfc/_565_ ( .A(\myfc/_316_ ), .Z(\src1 [5] ) );
BUF_X1 \myfc/_566_ ( .A(\EX_LS_result_reg [6] ), .Z(\myfc/_069_ ) );
BUF_X1 \myfc/_567_ ( .A(\src1_raw [6] ), .Z(\myfc/_221_ ) );
BUF_X1 \myfc/_568_ ( .A(\myfc/_317_ ), .Z(\src1 [6] ) );
BUF_X1 \myfc/_569_ ( .A(\EX_LS_result_reg [7] ), .Z(\myfc/_070_ ) );
BUF_X1 \myfc/_570_ ( .A(\src1_raw [7] ), .Z(\myfc/_222_ ) );
BUF_X1 \myfc/_571_ ( .A(\myfc/_318_ ), .Z(\src1 [7] ) );
BUF_X1 \myfc/_572_ ( .A(\EX_LS_result_reg [8] ), .Z(\myfc/_071_ ) );
BUF_X1 \myfc/_573_ ( .A(\src1_raw [8] ), .Z(\myfc/_223_ ) );
BUF_X1 \myfc/_574_ ( .A(\myfc/_319_ ), .Z(\src1 [8] ) );
BUF_X1 \myfc/_575_ ( .A(\EX_LS_result_reg [9] ), .Z(\myfc/_072_ ) );
BUF_X1 \myfc/_576_ ( .A(\src1_raw [9] ), .Z(\myfc/_224_ ) );
BUF_X1 \myfc/_577_ ( .A(\myfc/_320_ ), .Z(\src1 [9] ) );
BUF_X1 \myfc/_578_ ( .A(\EX_LS_result_reg [10] ), .Z(\myfc/_042_ ) );
BUF_X1 \myfc/_579_ ( .A(\src1_raw [10] ), .Z(\myfc/_194_ ) );
BUF_X1 \myfc/_580_ ( .A(\myfc/_290_ ), .Z(\src1 [10] ) );
BUF_X1 \myfc/_581_ ( .A(\EX_LS_result_reg [11] ), .Z(\myfc/_043_ ) );
BUF_X1 \myfc/_582_ ( .A(\src1_raw [11] ), .Z(\myfc/_195_ ) );
BUF_X1 \myfc/_583_ ( .A(\myfc/_291_ ), .Z(\src1 [11] ) );
BUF_X1 \myfc/_584_ ( .A(\EX_LS_result_reg [12] ), .Z(\myfc/_044_ ) );
BUF_X1 \myfc/_585_ ( .A(\src1_raw [12] ), .Z(\myfc/_196_ ) );
BUF_X1 \myfc/_586_ ( .A(\myfc/_292_ ), .Z(\src1 [12] ) );
BUF_X1 \myfc/_587_ ( .A(\EX_LS_result_reg [13] ), .Z(\myfc/_045_ ) );
BUF_X1 \myfc/_588_ ( .A(\src1_raw [13] ), .Z(\myfc/_197_ ) );
BUF_X1 \myfc/_589_ ( .A(\myfc/_293_ ), .Z(\src1 [13] ) );
BUF_X1 \myfc/_590_ ( .A(\EX_LS_result_reg [14] ), .Z(\myfc/_046_ ) );
BUF_X1 \myfc/_591_ ( .A(\src1_raw [14] ), .Z(\myfc/_198_ ) );
BUF_X1 \myfc/_592_ ( .A(\myfc/_294_ ), .Z(\src1 [14] ) );
BUF_X1 \myfc/_593_ ( .A(\EX_LS_result_reg [15] ), .Z(\myfc/_047_ ) );
BUF_X1 \myfc/_594_ ( .A(\src1_raw [15] ), .Z(\myfc/_199_ ) );
BUF_X1 \myfc/_595_ ( .A(\myfc/_295_ ), .Z(\src1 [15] ) );
BUF_X1 \myfc/_596_ ( .A(\EX_LS_result_reg [16] ), .Z(\myfc/_048_ ) );
BUF_X1 \myfc/_597_ ( .A(\src1_raw [16] ), .Z(\myfc/_200_ ) );
BUF_X1 \myfc/_598_ ( .A(\myfc/_296_ ), .Z(\src1 [16] ) );
BUF_X1 \myfc/_599_ ( .A(\EX_LS_result_reg [17] ), .Z(\myfc/_049_ ) );
BUF_X1 \myfc/_600_ ( .A(\src1_raw [17] ), .Z(\myfc/_201_ ) );
BUF_X1 \myfc/_601_ ( .A(\myfc/_297_ ), .Z(\src1 [17] ) );
BUF_X1 \myfc/_602_ ( .A(\EX_LS_result_reg [18] ), .Z(\myfc/_050_ ) );
BUF_X1 \myfc/_603_ ( .A(\src1_raw [18] ), .Z(\myfc/_202_ ) );
BUF_X1 \myfc/_604_ ( .A(\myfc/_298_ ), .Z(\src1 [18] ) );
BUF_X1 \myfc/_605_ ( .A(\EX_LS_result_reg [19] ), .Z(\myfc/_051_ ) );
BUF_X1 \myfc/_606_ ( .A(\src1_raw [19] ), .Z(\myfc/_203_ ) );
BUF_X1 \myfc/_607_ ( .A(\myfc/_299_ ), .Z(\src1 [19] ) );
BUF_X1 \myfc/_608_ ( .A(\EX_LS_result_reg [20] ), .Z(\myfc/_053_ ) );
BUF_X1 \myfc/_609_ ( .A(\src1_raw [20] ), .Z(\myfc/_205_ ) );
BUF_X1 \myfc/_610_ ( .A(\myfc/_301_ ), .Z(\src1 [20] ) );
BUF_X1 \myfc/_611_ ( .A(\EX_LS_result_reg [21] ), .Z(\myfc/_054_ ) );
BUF_X1 \myfc/_612_ ( .A(\src1_raw [21] ), .Z(\myfc/_206_ ) );
BUF_X1 \myfc/_613_ ( .A(\myfc/_302_ ), .Z(\src1 [21] ) );
BUF_X1 \myfc/_614_ ( .A(\EX_LS_result_reg [22] ), .Z(\myfc/_055_ ) );
BUF_X1 \myfc/_615_ ( .A(\src1_raw [22] ), .Z(\myfc/_207_ ) );
BUF_X1 \myfc/_616_ ( .A(\myfc/_303_ ), .Z(\src1 [22] ) );
BUF_X1 \myfc/_617_ ( .A(\EX_LS_result_reg [23] ), .Z(\myfc/_056_ ) );
BUF_X1 \myfc/_618_ ( .A(\src1_raw [23] ), .Z(\myfc/_208_ ) );
BUF_X1 \myfc/_619_ ( .A(\myfc/_304_ ), .Z(\src1 [23] ) );
BUF_X1 \myfc/_620_ ( .A(\EX_LS_result_reg [24] ), .Z(\myfc/_057_ ) );
BUF_X1 \myfc/_621_ ( .A(\src1_raw [24] ), .Z(\myfc/_209_ ) );
BUF_X1 \myfc/_622_ ( .A(\myfc/_305_ ), .Z(\src1 [24] ) );
BUF_X1 \myfc/_623_ ( .A(\EX_LS_result_reg [25] ), .Z(\myfc/_058_ ) );
BUF_X1 \myfc/_624_ ( .A(\src1_raw [25] ), .Z(\myfc/_210_ ) );
BUF_X1 \myfc/_625_ ( .A(\myfc/_306_ ), .Z(\src1 [25] ) );
BUF_X1 \myfc/_626_ ( .A(\EX_LS_result_reg [26] ), .Z(\myfc/_059_ ) );
BUF_X1 \myfc/_627_ ( .A(\src1_raw [26] ), .Z(\myfc/_211_ ) );
BUF_X1 \myfc/_628_ ( .A(\myfc/_307_ ), .Z(\src1 [26] ) );
BUF_X1 \myfc/_629_ ( .A(\EX_LS_result_reg [27] ), .Z(\myfc/_060_ ) );
BUF_X1 \myfc/_630_ ( .A(\src1_raw [27] ), .Z(\myfc/_212_ ) );
BUF_X1 \myfc/_631_ ( .A(\myfc/_308_ ), .Z(\src1 [27] ) );
BUF_X1 \myfc/_632_ ( .A(\EX_LS_result_reg [28] ), .Z(\myfc/_061_ ) );
BUF_X1 \myfc/_633_ ( .A(\src1_raw [28] ), .Z(\myfc/_213_ ) );
BUF_X1 \myfc/_634_ ( .A(\myfc/_309_ ), .Z(\src1 [28] ) );
BUF_X1 \myfc/_635_ ( .A(\EX_LS_result_reg [29] ), .Z(\myfc/_062_ ) );
BUF_X1 \myfc/_636_ ( .A(\src1_raw [29] ), .Z(\myfc/_214_ ) );
BUF_X1 \myfc/_637_ ( .A(\myfc/_310_ ), .Z(\src1 [29] ) );
BUF_X1 \myfc/_638_ ( .A(\EX_LS_result_reg [30] ), .Z(\myfc/_064_ ) );
BUF_X1 \myfc/_639_ ( .A(\src1_raw [30] ), .Z(\myfc/_216_ ) );
BUF_X1 \myfc/_640_ ( .A(\myfc/_312_ ), .Z(\src1 [30] ) );
BUF_X1 \myfc/_641_ ( .A(\EX_LS_result_reg [31] ), .Z(\myfc/_065_ ) );
BUF_X1 \myfc/_642_ ( .A(\src1_raw [31] ), .Z(\myfc/_217_ ) );
BUF_X1 \myfc/_643_ ( .A(\myfc/_313_ ), .Z(\src1 [31] ) );
BUF_X1 \myfc/_644_ ( .A(\ID_EX_rs2 [0] ), .Z(\myfc/_036_ ) );
BUF_X1 \myfc/_645_ ( .A(\ID_EX_rs2 [1] ), .Z(\myfc/_037_ ) );
BUF_X1 \myfc/_646_ ( .A(\ID_EX_rs2 [2] ), .Z(\myfc/_038_ ) );
BUF_X1 \myfc/_647_ ( .A(\ID_EX_rs2 [3] ), .Z(\myfc/_039_ ) );
BUF_X1 \myfc/_648_ ( .A(\ID_EX_rs2 [4] ), .Z(\myfc/_040_ ) );
BUF_X1 \myfc/_649_ ( .A(\EX_LS_result_reg [0] ), .Z(\myfc/_073_ ) );
BUF_X1 \myfc/_650_ ( .A(\src2_raw [0] ), .Z(\myfc/_225_ ) );
BUF_X1 \myfc/_651_ ( .A(\myfc/_321_ ), .Z(\src2 [0] ) );
BUF_X1 \myfc/_652_ ( .A(\EX_LS_result_reg [1] ), .Z(\myfc/_084_ ) );
BUF_X1 \myfc/_653_ ( .A(\src2_raw [1] ), .Z(\myfc/_236_ ) );
BUF_X1 \myfc/_654_ ( .A(\myfc/_332_ ), .Z(\src2 [1] ) );
BUF_X1 \myfc/_655_ ( .A(\EX_LS_result_reg [2] ), .Z(\myfc/_095_ ) );
BUF_X1 \myfc/_656_ ( .A(\src2_raw [2] ), .Z(\myfc/_247_ ) );
BUF_X1 \myfc/_657_ ( .A(\myfc/_343_ ), .Z(\src2 [2] ) );
BUF_X1 \myfc/_658_ ( .A(\EX_LS_result_reg [3] ), .Z(\myfc/_098_ ) );
BUF_X1 \myfc/_659_ ( .A(\src2_raw [3] ), .Z(\myfc/_250_ ) );
BUF_X1 \myfc/_660_ ( .A(\myfc/_346_ ), .Z(\src2 [3] ) );
BUF_X1 \myfc/_661_ ( .A(\EX_LS_result_reg [4] ), .Z(\myfc/_099_ ) );
BUF_X1 \myfc/_662_ ( .A(\src2_raw [4] ), .Z(\myfc/_251_ ) );
BUF_X1 \myfc/_663_ ( .A(\myfc/_347_ ), .Z(\src2 [4] ) );
BUF_X1 \myfc/_664_ ( .A(\EX_LS_result_reg [5] ), .Z(\myfc/_100_ ) );
BUF_X1 \myfc/_665_ ( .A(\src2_raw [5] ), .Z(\myfc/_252_ ) );
BUF_X1 \myfc/_666_ ( .A(\myfc/_348_ ), .Z(\src2 [5] ) );
BUF_X1 \myfc/_667_ ( .A(\EX_LS_result_reg [6] ), .Z(\myfc/_101_ ) );
BUF_X1 \myfc/_668_ ( .A(\src2_raw [6] ), .Z(\myfc/_253_ ) );
BUF_X1 \myfc/_669_ ( .A(\myfc/_349_ ), .Z(\src2 [6] ) );
BUF_X1 \myfc/_670_ ( .A(\EX_LS_result_reg [7] ), .Z(\myfc/_102_ ) );
BUF_X1 \myfc/_671_ ( .A(\src2_raw [7] ), .Z(\myfc/_254_ ) );
BUF_X1 \myfc/_672_ ( .A(\myfc/_350_ ), .Z(\src2 [7] ) );
BUF_X1 \myfc/_673_ ( .A(\EX_LS_result_reg [8] ), .Z(\myfc/_103_ ) );
BUF_X1 \myfc/_674_ ( .A(\src2_raw [8] ), .Z(\myfc/_255_ ) );
BUF_X1 \myfc/_675_ ( .A(\myfc/_351_ ), .Z(\src2 [8] ) );
BUF_X1 \myfc/_676_ ( .A(\EX_LS_result_reg [9] ), .Z(\myfc/_104_ ) );
BUF_X1 \myfc/_677_ ( .A(\src2_raw [9] ), .Z(\myfc/_256_ ) );
BUF_X1 \myfc/_678_ ( .A(\myfc/_352_ ), .Z(\src2 [9] ) );
BUF_X1 \myfc/_679_ ( .A(\EX_LS_result_reg [10] ), .Z(\myfc/_074_ ) );
BUF_X1 \myfc/_680_ ( .A(\src2_raw [10] ), .Z(\myfc/_226_ ) );
BUF_X1 \myfc/_681_ ( .A(\myfc/_322_ ), .Z(\src2 [10] ) );
BUF_X1 \myfc/_682_ ( .A(\EX_LS_result_reg [11] ), .Z(\myfc/_075_ ) );
BUF_X1 \myfc/_683_ ( .A(\src2_raw [11] ), .Z(\myfc/_227_ ) );
BUF_X1 \myfc/_684_ ( .A(\myfc/_323_ ), .Z(\src2 [11] ) );
BUF_X1 \myfc/_685_ ( .A(\EX_LS_result_reg [12] ), .Z(\myfc/_076_ ) );
BUF_X1 \myfc/_686_ ( .A(\src2_raw [12] ), .Z(\myfc/_228_ ) );
BUF_X1 \myfc/_687_ ( .A(\myfc/_324_ ), .Z(\src2 [12] ) );
BUF_X1 \myfc/_688_ ( .A(\EX_LS_result_reg [13] ), .Z(\myfc/_077_ ) );
BUF_X1 \myfc/_689_ ( .A(\src2_raw [13] ), .Z(\myfc/_229_ ) );
BUF_X1 \myfc/_690_ ( .A(\myfc/_325_ ), .Z(\src2 [13] ) );
BUF_X1 \myfc/_691_ ( .A(\EX_LS_result_reg [14] ), .Z(\myfc/_078_ ) );
BUF_X1 \myfc/_692_ ( .A(\src2_raw [14] ), .Z(\myfc/_230_ ) );
BUF_X1 \myfc/_693_ ( .A(\myfc/_326_ ), .Z(\src2 [14] ) );
BUF_X1 \myfc/_694_ ( .A(\EX_LS_result_reg [15] ), .Z(\myfc/_079_ ) );
BUF_X1 \myfc/_695_ ( .A(\src2_raw [15] ), .Z(\myfc/_231_ ) );
BUF_X1 \myfc/_696_ ( .A(\myfc/_327_ ), .Z(\src2 [15] ) );
BUF_X1 \myfc/_697_ ( .A(\EX_LS_result_reg [16] ), .Z(\myfc/_080_ ) );
BUF_X1 \myfc/_698_ ( .A(\src2_raw [16] ), .Z(\myfc/_232_ ) );
BUF_X1 \myfc/_699_ ( .A(\myfc/_328_ ), .Z(\src2 [16] ) );
BUF_X1 \myfc/_700_ ( .A(\EX_LS_result_reg [17] ), .Z(\myfc/_081_ ) );
BUF_X1 \myfc/_701_ ( .A(\src2_raw [17] ), .Z(\myfc/_233_ ) );
BUF_X1 \myfc/_702_ ( .A(\myfc/_329_ ), .Z(\src2 [17] ) );
BUF_X1 \myfc/_703_ ( .A(\EX_LS_result_reg [18] ), .Z(\myfc/_082_ ) );
BUF_X1 \myfc/_704_ ( .A(\src2_raw [18] ), .Z(\myfc/_234_ ) );
BUF_X1 \myfc/_705_ ( .A(\myfc/_330_ ), .Z(\src2 [18] ) );
BUF_X1 \myfc/_706_ ( .A(\EX_LS_result_reg [19] ), .Z(\myfc/_083_ ) );
BUF_X1 \myfc/_707_ ( .A(\src2_raw [19] ), .Z(\myfc/_235_ ) );
BUF_X1 \myfc/_708_ ( .A(\myfc/_331_ ), .Z(\src2 [19] ) );
BUF_X1 \myfc/_709_ ( .A(\EX_LS_result_reg [20] ), .Z(\myfc/_085_ ) );
BUF_X1 \myfc/_710_ ( .A(\src2_raw [20] ), .Z(\myfc/_237_ ) );
BUF_X1 \myfc/_711_ ( .A(\myfc/_333_ ), .Z(\src2 [20] ) );
BUF_X1 \myfc/_712_ ( .A(\EX_LS_result_reg [21] ), .Z(\myfc/_086_ ) );
BUF_X1 \myfc/_713_ ( .A(\src2_raw [21] ), .Z(\myfc/_238_ ) );
BUF_X1 \myfc/_714_ ( .A(\myfc/_334_ ), .Z(\src2 [21] ) );
BUF_X1 \myfc/_715_ ( .A(\EX_LS_result_reg [22] ), .Z(\myfc/_087_ ) );
BUF_X1 \myfc/_716_ ( .A(\src2_raw [22] ), .Z(\myfc/_239_ ) );
BUF_X1 \myfc/_717_ ( .A(\myfc/_335_ ), .Z(\src2 [22] ) );
BUF_X1 \myfc/_718_ ( .A(\EX_LS_result_reg [23] ), .Z(\myfc/_088_ ) );
BUF_X1 \myfc/_719_ ( .A(\src2_raw [23] ), .Z(\myfc/_240_ ) );
BUF_X1 \myfc/_720_ ( .A(\myfc/_336_ ), .Z(\src2 [23] ) );
BUF_X1 \myfc/_721_ ( .A(\EX_LS_result_reg [24] ), .Z(\myfc/_089_ ) );
BUF_X1 \myfc/_722_ ( .A(\src2_raw [24] ), .Z(\myfc/_241_ ) );
BUF_X1 \myfc/_723_ ( .A(\myfc/_337_ ), .Z(\src2 [24] ) );
BUF_X1 \myfc/_724_ ( .A(\EX_LS_result_reg [25] ), .Z(\myfc/_090_ ) );
BUF_X1 \myfc/_725_ ( .A(\src2_raw [25] ), .Z(\myfc/_242_ ) );
BUF_X1 \myfc/_726_ ( .A(\myfc/_338_ ), .Z(\src2 [25] ) );
BUF_X1 \myfc/_727_ ( .A(\EX_LS_result_reg [26] ), .Z(\myfc/_091_ ) );
BUF_X1 \myfc/_728_ ( .A(\src2_raw [26] ), .Z(\myfc/_243_ ) );
BUF_X1 \myfc/_729_ ( .A(\myfc/_339_ ), .Z(\src2 [26] ) );
BUF_X1 \myfc/_730_ ( .A(\EX_LS_result_reg [27] ), .Z(\myfc/_092_ ) );
BUF_X1 \myfc/_731_ ( .A(\src2_raw [27] ), .Z(\myfc/_244_ ) );
BUF_X1 \myfc/_732_ ( .A(\myfc/_340_ ), .Z(\src2 [27] ) );
BUF_X1 \myfc/_733_ ( .A(\EX_LS_result_reg [28] ), .Z(\myfc/_093_ ) );
BUF_X1 \myfc/_734_ ( .A(\src2_raw [28] ), .Z(\myfc/_245_ ) );
BUF_X1 \myfc/_735_ ( .A(\myfc/_341_ ), .Z(\src2 [28] ) );
BUF_X1 \myfc/_736_ ( .A(\EX_LS_result_reg [29] ), .Z(\myfc/_094_ ) );
BUF_X1 \myfc/_737_ ( .A(\src2_raw [29] ), .Z(\myfc/_246_ ) );
BUF_X1 \myfc/_738_ ( .A(\myfc/_342_ ), .Z(\src2 [29] ) );
BUF_X1 \myfc/_739_ ( .A(\EX_LS_result_reg [30] ), .Z(\myfc/_096_ ) );
BUF_X1 \myfc/_740_ ( .A(\src2_raw [30] ), .Z(\myfc/_248_ ) );
BUF_X1 \myfc/_741_ ( .A(\myfc/_344_ ), .Z(\src2 [30] ) );
BUF_X1 \myfc/_742_ ( .A(\EX_LS_result_reg [31] ), .Z(\myfc/_097_ ) );
BUF_X1 \myfc/_743_ ( .A(\src2_raw [31] ), .Z(\myfc/_249_ ) );
BUF_X1 \myfc/_744_ ( .A(\myfc/_345_ ), .Z(\src2 [31] ) );
BUF_X1 \myfc/_745_ ( .A(\ID_EX_csr [0] ), .Z(\myfc/_019_ ) );
BUF_X1 \myfc/_746_ ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(\myfc/_002_ ) );
BUF_X1 \myfc/_747_ ( .A(\ID_EX_csr [1] ), .Z(\myfc/_022_ ) );
BUF_X1 \myfc/_748_ ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(\myfc/_005_ ) );
BUF_X1 \myfc/_749_ ( .A(\ID_EX_csr [2] ), .Z(\myfc/_023_ ) );
BUF_X1 \myfc/_750_ ( .A(\EX_LS_dest_csreg_mem [2] ), .Z(\myfc/_006_ ) );
BUF_X1 \myfc/_751_ ( .A(\ID_EX_csr [3] ), .Z(\myfc/_024_ ) );
BUF_X1 \myfc/_752_ ( .A(\EX_LS_dest_csreg_mem [3] ), .Z(\myfc/_007_ ) );
BUF_X1 \myfc/_753_ ( .A(\ID_EX_csr [4] ), .Z(\myfc/_025_ ) );
BUF_X1 \myfc/_754_ ( .A(\EX_LS_dest_csreg_mem [4] ), .Z(\myfc/_008_ ) );
BUF_X1 \myfc/_755_ ( .A(\ID_EX_csr [5] ), .Z(\myfc/_026_ ) );
BUF_X1 \myfc/_756_ ( .A(\EX_LS_dest_csreg_mem [5] ), .Z(\myfc/_009_ ) );
BUF_X1 \myfc/_757_ ( .A(\ID_EX_csr [6] ), .Z(\myfc/_027_ ) );
BUF_X1 \myfc/_758_ ( .A(\EX_LS_dest_csreg_mem [6] ), .Z(\myfc/_010_ ) );
BUF_X1 \myfc/_759_ ( .A(\ID_EX_csr [7] ), .Z(\myfc/_028_ ) );
BUF_X1 \myfc/_760_ ( .A(\EX_LS_dest_csreg_mem [7] ), .Z(\myfc/_011_ ) );
BUF_X1 \myfc/_761_ ( .A(\ID_EX_csr [8] ), .Z(\myfc/_029_ ) );
BUF_X1 \myfc/_762_ ( .A(\EX_LS_dest_csreg_mem [8] ), .Z(\myfc/_012_ ) );
BUF_X1 \myfc/_763_ ( .A(\ID_EX_csr [9] ), .Z(\myfc/_030_ ) );
BUF_X1 \myfc/_764_ ( .A(\EX_LS_dest_csreg_mem [9] ), .Z(\myfc/_013_ ) );
BUF_X1 \myfc/_765_ ( .A(\ID_EX_csr [10] ), .Z(\myfc/_020_ ) );
BUF_X1 \myfc/_766_ ( .A(\EX_LS_dest_csreg_mem [10] ), .Z(\myfc/_003_ ) );
BUF_X1 \myfc/_767_ ( .A(\ID_EX_csr [11] ), .Z(\myfc/_021_ ) );
BUF_X1 \myfc/_768_ ( .A(\EX_LS_dest_csreg_mem [11] ), .Z(\myfc/_004_ ) );
BUF_X1 \myfc/_769_ ( .A(EX_LS_CSRegWrite ), .Z(\myfc/_000_ ) );
BUF_X1 \myfc/_770_ ( .A(\EX_LS_result_csreg_mem [0] ), .Z(\myfc/_105_ ) );
BUF_X1 \myfc/_771_ ( .A(\srccs_raw [0] ), .Z(\myfc/_257_ ) );
BUF_X1 \myfc/_772_ ( .A(\myfc/_353_ ), .Z(\srccs [0] ) );
BUF_X1 \myfc/_773_ ( .A(\EX_LS_result_csreg_mem [1] ), .Z(\myfc/_116_ ) );
BUF_X1 \myfc/_774_ ( .A(\srccs_raw [1] ), .Z(\myfc/_268_ ) );
BUF_X1 \myfc/_775_ ( .A(\myfc/_364_ ), .Z(\srccs [1] ) );
BUF_X1 \myfc/_776_ ( .A(\EX_LS_result_csreg_mem [2] ), .Z(\myfc/_127_ ) );
BUF_X1 \myfc/_777_ ( .A(\srccs_raw [2] ), .Z(\myfc/_279_ ) );
BUF_X1 \myfc/_778_ ( .A(\myfc/_375_ ), .Z(\srccs [2] ) );
BUF_X1 \myfc/_779_ ( .A(\EX_LS_result_csreg_mem [3] ), .Z(\myfc/_130_ ) );
BUF_X1 \myfc/_780_ ( .A(\srccs_raw [3] ), .Z(\myfc/_282_ ) );
BUF_X1 \myfc/_781_ ( .A(\myfc/_378_ ), .Z(\srccs [3] ) );
BUF_X1 \myfc/_782_ ( .A(\EX_LS_result_csreg_mem [4] ), .Z(\myfc/_131_ ) );
BUF_X1 \myfc/_783_ ( .A(\srccs_raw [4] ), .Z(\myfc/_283_ ) );
BUF_X1 \myfc/_784_ ( .A(\myfc/_379_ ), .Z(\srccs [4] ) );
BUF_X1 \myfc/_785_ ( .A(\EX_LS_result_csreg_mem [5] ), .Z(\myfc/_132_ ) );
BUF_X1 \myfc/_786_ ( .A(\srccs_raw [5] ), .Z(\myfc/_284_ ) );
BUF_X1 \myfc/_787_ ( .A(\myfc/_380_ ), .Z(\srccs [5] ) );
BUF_X1 \myfc/_788_ ( .A(\EX_LS_result_csreg_mem [6] ), .Z(\myfc/_133_ ) );
BUF_X1 \myfc/_789_ ( .A(\srccs_raw [6] ), .Z(\myfc/_285_ ) );
BUF_X1 \myfc/_790_ ( .A(\myfc/_381_ ), .Z(\srccs [6] ) );
BUF_X1 \myfc/_791_ ( .A(\EX_LS_result_csreg_mem [7] ), .Z(\myfc/_134_ ) );
BUF_X1 \myfc/_792_ ( .A(\srccs_raw [7] ), .Z(\myfc/_286_ ) );
BUF_X1 \myfc/_793_ ( .A(\myfc/_382_ ), .Z(\srccs [7] ) );
BUF_X1 \myfc/_794_ ( .A(\EX_LS_result_csreg_mem [8] ), .Z(\myfc/_135_ ) );
BUF_X1 \myfc/_795_ ( .A(\srccs_raw [8] ), .Z(\myfc/_287_ ) );
BUF_X1 \myfc/_796_ ( .A(\myfc/_383_ ), .Z(\srccs [8] ) );
BUF_X1 \myfc/_797_ ( .A(\EX_LS_result_csreg_mem [9] ), .Z(\myfc/_136_ ) );
BUF_X1 \myfc/_798_ ( .A(\srccs_raw [9] ), .Z(\myfc/_288_ ) );
BUF_X1 \myfc/_799_ ( .A(\myfc/_384_ ), .Z(\srccs [9] ) );
BUF_X1 \myfc/_800_ ( .A(\EX_LS_result_csreg_mem [10] ), .Z(\myfc/_106_ ) );
BUF_X1 \myfc/_801_ ( .A(\srccs_raw [10] ), .Z(\myfc/_258_ ) );
BUF_X1 \myfc/_802_ ( .A(\myfc/_354_ ), .Z(\srccs [10] ) );
BUF_X1 \myfc/_803_ ( .A(\EX_LS_result_csreg_mem [11] ), .Z(\myfc/_107_ ) );
BUF_X1 \myfc/_804_ ( .A(\srccs_raw [11] ), .Z(\myfc/_259_ ) );
BUF_X1 \myfc/_805_ ( .A(\myfc/_355_ ), .Z(\srccs [11] ) );
BUF_X1 \myfc/_806_ ( .A(\EX_LS_result_csreg_mem [12] ), .Z(\myfc/_108_ ) );
BUF_X1 \myfc/_807_ ( .A(\srccs_raw [12] ), .Z(\myfc/_260_ ) );
BUF_X1 \myfc/_808_ ( .A(\myfc/_356_ ), .Z(\srccs [12] ) );
BUF_X1 \myfc/_809_ ( .A(\EX_LS_result_csreg_mem [13] ), .Z(\myfc/_109_ ) );
BUF_X1 \myfc/_810_ ( .A(\srccs_raw [13] ), .Z(\myfc/_261_ ) );
BUF_X1 \myfc/_811_ ( .A(\myfc/_357_ ), .Z(\srccs [13] ) );
BUF_X1 \myfc/_812_ ( .A(\EX_LS_result_csreg_mem [14] ), .Z(\myfc/_110_ ) );
BUF_X1 \myfc/_813_ ( .A(\srccs_raw [14] ), .Z(\myfc/_262_ ) );
BUF_X1 \myfc/_814_ ( .A(\myfc/_358_ ), .Z(\srccs [14] ) );
BUF_X1 \myfc/_815_ ( .A(\EX_LS_result_csreg_mem [15] ), .Z(\myfc/_111_ ) );
BUF_X1 \myfc/_816_ ( .A(\srccs_raw [15] ), .Z(\myfc/_263_ ) );
BUF_X1 \myfc/_817_ ( .A(\myfc/_359_ ), .Z(\srccs [15] ) );
BUF_X1 \myfc/_818_ ( .A(\EX_LS_result_csreg_mem [16] ), .Z(\myfc/_112_ ) );
BUF_X1 \myfc/_819_ ( .A(\srccs_raw [16] ), .Z(\myfc/_264_ ) );
BUF_X1 \myfc/_820_ ( .A(\myfc/_360_ ), .Z(\srccs [16] ) );
BUF_X1 \myfc/_821_ ( .A(\EX_LS_result_csreg_mem [17] ), .Z(\myfc/_113_ ) );
BUF_X1 \myfc/_822_ ( .A(\srccs_raw [17] ), .Z(\myfc/_265_ ) );
BUF_X1 \myfc/_823_ ( .A(\myfc/_361_ ), .Z(\srccs [17] ) );
BUF_X1 \myfc/_824_ ( .A(\EX_LS_result_csreg_mem [18] ), .Z(\myfc/_114_ ) );
BUF_X1 \myfc/_825_ ( .A(\srccs_raw [18] ), .Z(\myfc/_266_ ) );
BUF_X1 \myfc/_826_ ( .A(\myfc/_362_ ), .Z(\srccs [18] ) );
BUF_X1 \myfc/_827_ ( .A(\EX_LS_result_csreg_mem [19] ), .Z(\myfc/_115_ ) );
BUF_X1 \myfc/_828_ ( .A(\srccs_raw [19] ), .Z(\myfc/_267_ ) );
BUF_X1 \myfc/_829_ ( .A(\myfc/_363_ ), .Z(\srccs [19] ) );
BUF_X1 \myfc/_830_ ( .A(\EX_LS_result_csreg_mem [20] ), .Z(\myfc/_117_ ) );
BUF_X1 \myfc/_831_ ( .A(\srccs_raw [20] ), .Z(\myfc/_269_ ) );
BUF_X1 \myfc/_832_ ( .A(\myfc/_365_ ), .Z(\srccs [20] ) );
BUF_X1 \myfc/_833_ ( .A(\EX_LS_result_csreg_mem [21] ), .Z(\myfc/_118_ ) );
BUF_X1 \myfc/_834_ ( .A(\srccs_raw [21] ), .Z(\myfc/_270_ ) );
BUF_X1 \myfc/_835_ ( .A(\myfc/_366_ ), .Z(\srccs [21] ) );
BUF_X1 \myfc/_836_ ( .A(\EX_LS_result_csreg_mem [22] ), .Z(\myfc/_119_ ) );
BUF_X1 \myfc/_837_ ( .A(\srccs_raw [22] ), .Z(\myfc/_271_ ) );
BUF_X1 \myfc/_838_ ( .A(\myfc/_367_ ), .Z(\srccs [22] ) );
BUF_X1 \myfc/_839_ ( .A(\EX_LS_result_csreg_mem [23] ), .Z(\myfc/_120_ ) );
BUF_X1 \myfc/_840_ ( .A(\srccs_raw [23] ), .Z(\myfc/_272_ ) );
BUF_X1 \myfc/_841_ ( .A(\myfc/_368_ ), .Z(\srccs [23] ) );
BUF_X1 \myfc/_842_ ( .A(\EX_LS_result_csreg_mem [24] ), .Z(\myfc/_121_ ) );
BUF_X1 \myfc/_843_ ( .A(\srccs_raw [24] ), .Z(\myfc/_273_ ) );
BUF_X1 \myfc/_844_ ( .A(\myfc/_369_ ), .Z(\srccs [24] ) );
BUF_X1 \myfc/_845_ ( .A(\EX_LS_result_csreg_mem [25] ), .Z(\myfc/_122_ ) );
BUF_X1 \myfc/_846_ ( .A(\srccs_raw [25] ), .Z(\myfc/_274_ ) );
BUF_X1 \myfc/_847_ ( .A(\myfc/_370_ ), .Z(\srccs [25] ) );
BUF_X1 \myfc/_848_ ( .A(\EX_LS_result_csreg_mem [26] ), .Z(\myfc/_123_ ) );
BUF_X1 \myfc/_849_ ( .A(\srccs_raw [26] ), .Z(\myfc/_275_ ) );
BUF_X1 \myfc/_850_ ( .A(\myfc/_371_ ), .Z(\srccs [26] ) );
BUF_X1 \myfc/_851_ ( .A(\EX_LS_result_csreg_mem [27] ), .Z(\myfc/_124_ ) );
BUF_X1 \myfc/_852_ ( .A(\srccs_raw [27] ), .Z(\myfc/_276_ ) );
BUF_X1 \myfc/_853_ ( .A(\myfc/_372_ ), .Z(\srccs [27] ) );
BUF_X1 \myfc/_854_ ( .A(\EX_LS_result_csreg_mem [28] ), .Z(\myfc/_125_ ) );
BUF_X1 \myfc/_855_ ( .A(\srccs_raw [28] ), .Z(\myfc/_277_ ) );
BUF_X1 \myfc/_856_ ( .A(\myfc/_373_ ), .Z(\srccs [28] ) );
BUF_X1 \myfc/_857_ ( .A(\EX_LS_result_csreg_mem [29] ), .Z(\myfc/_126_ ) );
BUF_X1 \myfc/_858_ ( .A(\srccs_raw [29] ), .Z(\myfc/_278_ ) );
BUF_X1 \myfc/_859_ ( .A(\myfc/_374_ ), .Z(\srccs [29] ) );
BUF_X1 \myfc/_860_ ( .A(\EX_LS_result_csreg_mem [30] ), .Z(\myfc/_128_ ) );
BUF_X1 \myfc/_861_ ( .A(\srccs_raw [30] ), .Z(\myfc/_280_ ) );
BUF_X1 \myfc/_862_ ( .A(\myfc/_376_ ), .Z(\srccs [30] ) );
BUF_X1 \myfc/_863_ ( .A(\EX_LS_result_csreg_mem [31] ), .Z(\myfc/_129_ ) );
BUF_X1 \myfc/_864_ ( .A(\srccs_raw [31] ), .Z(\myfc/_281_ ) );
BUF_X1 \myfc/_865_ ( .A(\myfc/_377_ ), .Z(\srccs [31] ) );
INV_X1 \myidu/_1009_ ( .A(\myidu/_0802_ ), .ZN(\myidu/_0188_ ) );
NOR2_X1 \myidu/_1010_ ( .A1(\myidu/_0188_ ), .A2(\myidu/_0777_ ), .ZN(\myidu/_0189_ ) );
INV_X1 \myidu/_1011_ ( .A(\myidu/_0182_ ), .ZN(\myidu/_0190_ ) );
NOR2_X1 \myidu/_1012_ ( .A1(\myidu/_0190_ ), .A2(\myidu/_0181_ ), .ZN(\myidu/_0191_ ) );
INV_X1 \myidu/_1013_ ( .A(\myidu/_0183_ ), .ZN(\myidu/_0192_ ) );
NOR2_X1 \myidu/_1014_ ( .A1(\myidu/_0192_ ), .A2(\myidu/_0158_ ), .ZN(\myidu/_0193_ ) );
NOR2_X1 \myidu/_1015_ ( .A1(\myidu/_0160_ ), .A2(\myidu/_0159_ ), .ZN(\myidu/_0194_ ) );
AND3_X1 \myidu/_1016_ ( .A1(\myidu/_0191_ ), .A2(\myidu/_0193_ ), .A3(\myidu/_0194_ ), .ZN(\myidu/_0195_ ) );
AND3_X1 \myidu/_1017_ ( .A1(\myidu/_0166_ ), .A2(\myidu/_0155_ ), .A3(\myidu/_0177_ ), .ZN(\myidu/_0196_ ) );
INV_X1 \myidu/_1018_ ( .A(\myidu/_0180_ ), .ZN(\myidu/_0197_ ) );
AND2_X1 \myidu/_1019_ ( .A1(\myidu/_0196_ ), .A2(\myidu/_0197_ ), .ZN(\myidu/_0198_ ) );
AND2_X1 \myidu/_1020_ ( .A1(\myidu/_0195_ ), .A2(\myidu/_0198_ ), .ZN(\myidu/_0199_ ) );
INV_X16 \myidu/_1021_ ( .A(\myidu/_0158_ ), .ZN(\myidu/_0200_ ) );
NOR2_X4 \myidu/_1022_ ( .A1(\myidu/_0200_ ), .A2(\myidu/_0183_ ), .ZN(\myidu/_0201_ ) );
AND2_X4 \myidu/_1023_ ( .A1(\myidu/_0166_ ), .A2(\myidu/_0155_ ), .ZN(\myidu/_0202_ ) );
NOR2_X4 \myidu/_1024_ ( .A1(\myidu/_0180_ ), .A2(\myidu/_0177_ ), .ZN(\myidu/_0203_ ) );
AND3_X2 \myidu/_1025_ ( .A1(\myidu/_0201_ ), .A2(\myidu/_0202_ ), .A3(\myidu/_0203_ ), .ZN(\myidu/_0204_ ) );
INV_X1 \myidu/_1026_ ( .A(\myidu/_0181_ ), .ZN(\myidu/_0205_ ) );
NOR2_X1 \myidu/_1027_ ( .A1(\myidu/_0205_ ), .A2(\myidu/_0182_ ), .ZN(\myidu/_0206_ ) );
AND2_X4 \myidu/_1028_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0206_ ), .ZN(\myidu/_0207_ ) );
INV_X1 \myidu/_1029_ ( .A(\myidu/_0159_ ), .ZN(\myidu/_0208_ ) );
NOR2_X2 \myidu/_1030_ ( .A1(\myidu/_0208_ ), .A2(\myidu/_0160_ ), .ZN(\myidu/_0209_ ) );
AND2_X4 \myidu/_1031_ ( .A1(\myidu/_0207_ ), .A2(\myidu/_0209_ ), .ZN(\myidu/_0210_ ) );
AND2_X4 \myidu/_1032_ ( .A1(\myidu/_0202_ ), .A2(\myidu/_0203_ ), .ZN(\myidu/_0211_ ) );
NOR2_X1 \myidu/_1033_ ( .A1(\myidu/_0183_ ), .A2(\myidu/_0158_ ), .ZN(\myidu/_0212_ ) );
AND3_X1 \myidu/_1034_ ( .A1(\myidu/_0211_ ), .A2(\myidu/_0212_ ), .A3(\myidu/_0206_ ), .ZN(\myidu/_0213_ ) );
AOI211_X2 \myidu/_1035_ ( .A(\myidu/_0199_ ), .B(\myidu/_0210_ ), .C1(\myidu/_0209_ ), .C2(\myidu/_0213_ ), .ZN(\myidu/_0214_ ) );
NOR2_X1 \myidu/_1036_ ( .A1(\myidu/_0182_ ), .A2(\myidu/_0181_ ), .ZN(\myidu/_0215_ ) );
AND2_X1 \myidu/_1037_ ( .A1(\myidu/_0201_ ), .A2(\myidu/_0215_ ), .ZN(\myidu/_0216_ ) );
AND3_X1 \myidu/_1038_ ( .A1(\myidu/_0202_ ), .A2(\myidu/_0208_ ), .A3(\myidu/_0203_ ), .ZN(\myidu/_0217_ ) );
AND2_X1 \myidu/_1039_ ( .A1(\myidu/_0216_ ), .A2(\myidu/_0217_ ), .ZN(\myidu/_0218_ ) );
INV_X1 \myidu/_1040_ ( .A(\myidu/_0218_ ), .ZN(\myidu/_0219_ ) );
AND2_X2 \myidu/_1041_ ( .A1(\myidu/_0211_ ), .A2(\myidu/_0212_ ), .ZN(\myidu/_0220_ ) );
AND2_X2 \myidu/_1042_ ( .A1(\myidu/_0160_ ), .A2(\myidu/_0159_ ), .ZN(\myidu/_0221_ ) );
INV_X1 \myidu/_1043_ ( .A(\myidu/_0221_ ), .ZN(\myidu/_0222_ ) );
NAND3_X1 \myidu/_1044_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0222_ ), .A3(\myidu/_0215_ ), .ZN(\myidu/_0223_ ) );
AND3_X2 \myidu/_1045_ ( .A1(\myidu/_0214_ ), .A2(\myidu/_0219_ ), .A3(\myidu/_0223_ ), .ZN(\myidu/_0224_ ) );
NAND3_X1 \myidu/_1046_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0159_ ), .A3(\myidu/_0206_ ), .ZN(\myidu/_0225_ ) );
INV_X1 \myidu/_1047_ ( .A(\myidu/_0160_ ), .ZN(\myidu/_0226_ ) );
NOR2_X1 \myidu/_1048_ ( .A1(\myidu/_0225_ ), .A2(\myidu/_0226_ ), .ZN(\myidu/_0227_ ) );
INV_X1 \myidu/_1049_ ( .A(\myidu/_0209_ ), .ZN(\myidu/_0228_ ) );
AOI21_X1 \myidu/_1050_ ( .A(\myidu/_0227_ ), .B1(\myidu/_0228_ ), .B2(\myidu/_0213_ ), .ZN(\myidu/_0229_ ) );
AND2_X1 \myidu/_1051_ ( .A1(\myidu/_0224_ ), .A2(\myidu/_0229_ ), .ZN(\myidu/_0230_ ) );
AND4_X1 \myidu/_1052_ ( .A1(\myidu/_0182_ ), .A2(\myidu/_0200_ ), .A3(\myidu/_0181_ ), .A4(\myidu/_0183_ ), .ZN(\myidu/_0231_ ) );
AND2_X1 \myidu/_1053_ ( .A1(\myidu/_0211_ ), .A2(\myidu/_0231_ ), .ZN(\myidu/_0232_ ) );
AND2_X4 \myidu/_1054_ ( .A1(\myidu/_0232_ ), .A2(\myidu/_0159_ ), .ZN(\myidu/_0233_ ) );
AND4_X1 \myidu/_1055_ ( .A1(\myidu/_0182_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0183_ ), .A4(\myidu/_0158_ ), .ZN(\myidu/_0234_ ) );
AND2_X1 \myidu/_1056_ ( .A1(\myidu/_0211_ ), .A2(\myidu/_0234_ ), .ZN(\myidu/_0235_ ) );
NOR2_X4 \myidu/_1057_ ( .A1(\myidu/_0233_ ), .A2(\myidu/_0235_ ), .ZN(\myidu/_0236_ ) );
AND2_X2 \myidu/_1058_ ( .A1(\myidu/_0230_ ), .A2(\myidu/_0236_ ), .ZN(\myidu/_0237_ ) );
INV_X1 \myidu/_1059_ ( .A(\myidu/_0237_ ), .ZN(\myidu/_0238_ ) );
XNOR2_X1 \myidu/_1060_ ( .A(\myidu/_0162_ ), .B(\myidu/_0773_ ), .ZN(\myidu/_0239_ ) );
XNOR2_X1 \myidu/_1061_ ( .A(\myidu/_0164_ ), .B(\myidu/_0775_ ), .ZN(\myidu/_0240_ ) );
XNOR2_X1 \myidu/_1062_ ( .A(\myidu/_0161_ ), .B(\myidu/_0772_ ), .ZN(\myidu/_0241_ ) );
XNOR2_X1 \myidu/_1063_ ( .A(\myidu/_0163_ ), .B(\myidu/_0774_ ), .ZN(\myidu/_0242_ ) );
NAND4_X1 \myidu/_1064_ ( .A1(\myidu/_0239_ ), .A2(\myidu/_0240_ ), .A3(\myidu/_0241_ ), .A4(\myidu/_0242_ ), .ZN(\myidu/_0243_ ) );
XOR2_X1 \myidu/_1065_ ( .A(\myidu/_0165_ ), .B(\myidu/_0776_ ), .Z(\myidu/_0244_ ) );
NOR2_X1 \myidu/_1066_ ( .A1(\myidu/_0243_ ), .A2(\myidu/_0244_ ), .ZN(\myidu/_0245_ ) );
INV_X1 \myidu/_1067_ ( .A(\myidu/_0800_ ), .ZN(\myidu/_0246_ ) );
AND2_X1 \myidu/_1068_ ( .A1(\myidu/_0246_ ), .A2(\myidu/_0799_ ), .ZN(\myidu/_0247_ ) );
AND2_X1 \myidu/_1069_ ( .A1(\myidu/_0247_ ), .A2(\myidu/_0798_ ), .ZN(\myidu/_0248_ ) );
AND2_X1 \myidu/_1070_ ( .A1(\myidu/_0245_ ), .A2(\myidu/_0248_ ), .ZN(\myidu/_0249_ ) );
NAND2_X1 \myidu/_1071_ ( .A1(\myidu/_0238_ ), .A2(\myidu/_0249_ ), .ZN(\myidu/_0250_ ) );
XNOR2_X1 \myidu/_1072_ ( .A(\myidu/_0776_ ), .B(\myidu/_0171_ ), .ZN(\myidu/_0251_ ) );
XNOR2_X1 \myidu/_1073_ ( .A(\myidu/_0775_ ), .B(\myidu/_0170_ ), .ZN(\myidu/_0252_ ) );
XNOR2_X1 \myidu/_1074_ ( .A(\myidu/_0772_ ), .B(\myidu/_0167_ ), .ZN(\myidu/_0253_ ) );
NAND4_X1 \myidu/_1075_ ( .A1(\myidu/_0248_ ), .A2(\myidu/_0251_ ), .A3(\myidu/_0252_ ), .A4(\myidu/_0253_ ), .ZN(\myidu/_0254_ ) );
XOR2_X1 \myidu/_1076_ ( .A(\myidu/_0773_ ), .B(\myidu/_0168_ ), .Z(\myidu/_0255_ ) );
XOR2_X1 \myidu/_1077_ ( .A(\myidu/_0774_ ), .B(\myidu/_0169_ ), .Z(\myidu/_0256_ ) );
NOR3_X1 \myidu/_1078_ ( .A1(\myidu/_0254_ ), .A2(\myidu/_0255_ ), .A3(\myidu/_0256_ ), .ZN(\myidu/_0257_ ) );
OR2_X1 \myidu/_1079_ ( .A1(\myidu/_0249_ ), .A2(\myidu/_0257_ ), .ZN(\myidu/_0258_ ) );
AND3_X2 \myidu/_1080_ ( .A1(\myidu/_0211_ ), .A2(\myidu/_0194_ ), .A3(\myidu/_0191_ ), .ZN(\myidu/_0259_ ) );
AND2_X2 \myidu/_1081_ ( .A1(\myidu/_0259_ ), .A2(\myidu/_0192_ ), .ZN(\myidu/_0260_ ) );
INV_X1 \myidu/_1082_ ( .A(\myidu/_0260_ ), .ZN(\myidu/_0261_ ) );
NAND3_X1 \myidu/_1083_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0209_ ), .A3(\myidu/_0191_ ), .ZN(\myidu/_0262_ ) );
NAND2_X4 \myidu/_1084_ ( .A1(\myidu/_0261_ ), .A2(\myidu/_0262_ ), .ZN(\myidu/_0263_ ) );
AND3_X1 \myidu/_1085_ ( .A1(\myidu/_0205_ ), .A2(\myidu/_0182_ ), .A3(\myidu/_0160_ ), .ZN(\myidu/_0264_ ) );
AND2_X4 \myidu/_1086_ ( .A1(\myidu/_0211_ ), .A2(\myidu/_0264_ ), .ZN(\myidu/_0265_ ) );
OR2_X4 \myidu/_1087_ ( .A1(\myidu/_0259_ ), .A2(\myidu/_0265_ ), .ZN(\myidu/_0266_ ) );
AND2_X4 \myidu/_1088_ ( .A1(\myidu/_0266_ ), .A2(\myidu/_0183_ ), .ZN(\myidu/_0267_ ) );
NOR2_X4 \myidu/_1089_ ( .A1(\myidu/_0263_ ), .A2(\myidu/_0267_ ), .ZN(\myidu/_0268_ ) );
NOR2_X1 \myidu/_1090_ ( .A1(\myidu/_0172_ ), .A2(\myidu/_0173_ ), .ZN(\myidu/_0269_ ) );
AND3_X1 \myidu/_1091_ ( .A1(\myidu/_0269_ ), .A2(\myidu/_0160_ ), .A3(\myidu/_0208_ ), .ZN(\myidu/_0270_ ) );
NOR2_X1 \myidu/_1092_ ( .A1(\myidu/_0176_ ), .A2(\myidu/_0175_ ), .ZN(\myidu/_0271_ ) );
INV_X1 \myidu/_1093_ ( .A(\myidu/_0174_ ), .ZN(\myidu/_0272_ ) );
AND3_X1 \myidu/_1094_ ( .A1(\myidu/_0271_ ), .A2(\myidu/_0272_ ), .A3(\myidu/_0178_ ), .ZN(\myidu/_0273_ ) );
NOR2_X1 \myidu/_1095_ ( .A1(\myidu/_0174_ ), .A2(\myidu/_0178_ ), .ZN(\myidu/_0274_ ) );
AND2_X1 \myidu/_1096_ ( .A1(\myidu/_0271_ ), .A2(\myidu/_0274_ ), .ZN(\myidu/_0275_ ) );
OAI21_X1 \myidu/_1097_ ( .A(\myidu/_0270_ ), .B1(\myidu/_0273_ ), .B2(\myidu/_0275_ ), .ZN(\myidu/_0276_ ) );
INV_X1 \myidu/_1098_ ( .A(\myidu/_0276_ ), .ZN(\myidu/_0277_ ) );
INV_X1 \myidu/_1099_ ( .A(\myidu/_0179_ ), .ZN(\myidu/_0278_ ) );
AND3_X2 \myidu/_1100_ ( .A1(\myidu/_0278_ ), .A2(\myidu/_0182_ ), .A3(\myidu/_0181_ ), .ZN(\myidu/_0279_ ) );
AND2_X1 \myidu/_1101_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0279_ ), .ZN(\myidu/_0280_ ) );
NAND2_X1 \myidu/_1102_ ( .A1(\myidu/_0277_ ), .A2(\myidu/_0280_ ), .ZN(\myidu/_0281_ ) );
INV_X1 \myidu/_1103_ ( .A(\myidu/_0172_ ), .ZN(\myidu/_0282_ ) );
INV_X1 \myidu/_1104_ ( .A(\myidu/_0173_ ), .ZN(\myidu/_0283_ ) );
AND4_X1 \myidu/_1105_ ( .A1(\myidu/_0226_ ), .A2(\myidu/_0282_ ), .A3(\myidu/_0283_ ), .A4(\myidu/_0159_ ), .ZN(\myidu/_0284_ ) );
AND2_X1 \myidu/_1106_ ( .A1(\myidu/_0275_ ), .A2(\myidu/_0284_ ), .ZN(\myidu/_0285_ ) );
NAND3_X1 \myidu/_1107_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0285_ ), .A3(\myidu/_0279_ ), .ZN(\myidu/_0286_ ) );
AND2_X1 \myidu/_1108_ ( .A1(\myidu/_0269_ ), .A2(\myidu/_0194_ ), .ZN(\myidu/_0287_ ) );
NAND4_X1 \myidu/_1109_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0279_ ), .A3(\myidu/_0273_ ), .A4(\myidu/_0287_ ), .ZN(\myidu/_0288_ ) );
AND3_X1 \myidu/_1110_ ( .A1(\myidu/_0281_ ), .A2(\myidu/_0286_ ), .A3(\myidu/_0288_ ), .ZN(\myidu/_0289_ ) );
BUF_X4 \myidu/_1111_ ( .A(\myidu/_0278_ ), .Z(\myidu/_0290_ ) );
AND3_X1 \myidu/_1112_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0290_ ), .A3(\myidu/_0206_ ), .ZN(\myidu/_0291_ ) );
AND2_X1 \myidu/_1113_ ( .A1(\myidu/_0291_ ), .A2(\myidu/_0277_ ), .ZN(\myidu/_0292_ ) );
AND2_X2 \myidu/_1114_ ( .A1(\myidu/_0275_ ), .A2(\myidu/_0287_ ), .ZN(\myidu/_0293_ ) );
AND2_X1 \myidu/_1115_ ( .A1(\myidu/_0291_ ), .A2(\myidu/_0293_ ), .ZN(\myidu/_0294_ ) );
NOR2_X1 \myidu/_1116_ ( .A1(\myidu/_0292_ ), .A2(\myidu/_0294_ ), .ZN(\myidu/_0295_ ) );
NAND3_X1 \myidu/_1117_ ( .A1(\myidu/_0268_ ), .A2(\myidu/_0289_ ), .A3(\myidu/_0295_ ), .ZN(\myidu/_0296_ ) );
CLKBUF_X2 \myidu/_1118_ ( .A(\myidu/_0211_ ), .Z(\myidu/_0297_ ) );
AND3_X1 \myidu/_1119_ ( .A1(\myidu/_0221_ ), .A2(\myidu/_0271_ ), .A3(\myidu/_0274_ ), .ZN(\myidu/_0298_ ) );
AND2_X1 \myidu/_1120_ ( .A1(\myidu/_0298_ ), .A2(\myidu/_0269_ ), .ZN(\myidu/_0299_ ) );
AND2_X1 \myidu/_1121_ ( .A1(\myidu/_0182_ ), .A2(\myidu/_0181_ ), .ZN(\myidu/_0300_ ) );
BUF_X2 \myidu/_1122_ ( .A(\myidu/_0300_ ), .Z(\myidu/_0301_ ) );
CLKBUF_X2 \myidu/_1123_ ( .A(\myidu/_0301_ ), .Z(\myidu/_0302_ ) );
CLKBUF_X2 \myidu/_1124_ ( .A(\myidu/_0212_ ), .Z(\myidu/_0303_ ) );
AND4_X1 \myidu/_1125_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0299_ ), .A3(\myidu/_0302_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0304_ ) );
AND2_X1 \myidu/_1126_ ( .A1(\myidu/_0270_ ), .A2(\myidu/_0275_ ), .ZN(\myidu/_0305_ ) );
AND4_X1 \myidu/_1127_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0305_ ), .A3(\myidu/_0301_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0306_ ) );
OAI21_X1 \myidu/_1128_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0304_ ), .B2(\myidu/_0306_ ), .ZN(\myidu/_0307_ ) );
CLKBUF_X2 \myidu/_1129_ ( .A(\myidu/_0201_ ), .Z(\myidu/_0308_ ) );
AND4_X1 \myidu/_1130_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0299_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0302_ ), .ZN(\myidu/_0309_ ) );
AND4_X1 \myidu/_1131_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0293_ ), .A3(\myidu/_0302_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0310_ ) );
OAI21_X1 \myidu/_1132_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0309_ ), .B2(\myidu/_0310_ ), .ZN(\myidu/_0311_ ) );
AND4_X1 \myidu/_1133_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0293_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0302_ ), .ZN(\myidu/_0312_ ) );
AND4_X1 \myidu/_1134_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0285_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0302_ ), .ZN(\myidu/_0313_ ) );
OAI21_X1 \myidu/_1135_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0312_ ), .B2(\myidu/_0313_ ), .ZN(\myidu/_0314_ ) );
NAND3_X1 \myidu/_1136_ ( .A1(\myidu/_0307_ ), .A2(\myidu/_0311_ ), .A3(\myidu/_0314_ ), .ZN(\myidu/_0315_ ) );
OAI21_X1 \myidu/_1137_ ( .A(\myidu/_0258_ ), .B1(\myidu/_0296_ ), .B2(\myidu/_0315_ ), .ZN(\myidu/_0316_ ) );
NAND2_X1 \myidu/_1138_ ( .A1(\myidu/_0250_ ), .A2(\myidu/_0316_ ), .ZN(\myidu/_0317_ ) );
INV_X1 \myidu/_1139_ ( .A(\myidu/_0317_ ), .ZN(\myidu/_0318_ ) );
AND2_X1 \myidu/_1140_ ( .A1(\myidu/_0778_ ), .A2(\myidu/_0801_ ), .ZN(\myidu/_0319_ ) );
BUF_X4 \myidu/_1141_ ( .A(\myidu/_0319_ ), .Z(\myidu/_0320_ ) );
AOI221_X4 \myidu/_1142_ ( .A(\myidu/_0189_ ), .B1(\myidu/_0187_ ), .B2(\myidu/_0792_ ), .C1(\myidu/_0318_ ), .C2(\myidu/_0320_ ), .ZN(\myidu/_0321_ ) );
NOR2_X1 \myidu/_1143_ ( .A1(\myidu/_0321_ ), .A2(\myidu/_0789_ ), .ZN(\myidu/_0005_ ) );
INV_X1 \myidu/_1144_ ( .A(\myidu/_0789_ ), .ZN(\myidu/_0322_ ) );
BUF_X4 \myidu/_1145_ ( .A(\myidu/_0322_ ), .Z(\myidu/_0323_ ) );
NAND3_X1 \myidu/_1146_ ( .A1(\myidu/_0323_ ), .A2(\myidu/_0777_ ), .A3(\myidu/_0802_ ), .ZN(\myidu/_0324_ ) );
BUF_X4 \myidu/_1147_ ( .A(\myidu/_0323_ ), .Z(\myidu/_0325_ ) );
INV_X1 \myidu/_1148_ ( .A(\myidu/_0778_ ), .ZN(\myidu/_0326_ ) );
OAI211_X2 \myidu/_1149_ ( .A(\myidu/_0324_ ), .B(\myidu/_0325_ ), .C1(\myidu/_0326_ ), .C2(\myidu/_0801_ ), .ZN(\myidu/_0004_ ) );
INV_X1 \myidu/_1150_ ( .A(\myidu/_0316_ ), .ZN(\myidu/_0327_ ) );
NAND4_X1 \myidu/_1151_ ( .A1(\myidu/_0327_ ), .A2(\myidu/_0778_ ), .A3(\myidu/_0323_ ), .A4(\myidu/_0801_ ), .ZN(\myidu/_0328_ ) );
INV_X1 \myidu/_1152_ ( .A(\myidu/_0792_ ), .ZN(\myidu/_0329_ ) );
OR3_X1 \myidu/_1153_ ( .A1(\myidu/_0329_ ), .A2(\myidu/_0789_ ), .A3(\myidu/_0187_ ), .ZN(\myidu/_0330_ ) );
NAND4_X1 \myidu/_1154_ ( .A1(\myidu/_0238_ ), .A2(\myidu/_0323_ ), .A3(\myidu/_0801_ ), .A4(\myidu/_0249_ ), .ZN(\myidu/_0331_ ) );
OAI211_X2 \myidu/_1155_ ( .A(\myidu/_0328_ ), .B(\myidu/_0330_ ), .C1(\myidu/_0326_ ), .C2(\myidu/_0331_ ), .ZN(\myidu/_0006_ ) );
INV_X1 \myidu/_1156_ ( .A(\myidu/_0236_ ), .ZN(\myidu/_0332_ ) );
BUF_X2 \myidu/_1157_ ( .A(\myidu/_0332_ ), .Z(\myidu/_0333_ ) );
AOI22_X1 \myidu/_1158_ ( .A1(\myidu/_0184_ ), .A2(\myidu/_0263_ ), .B1(\myidu/_0333_ ), .B2(\myidu/_0161_ ), .ZN(\myidu/_0334_ ) );
INV_X1 \myidu/_1159_ ( .A(\myidu/_0230_ ), .ZN(\myidu/_0335_ ) );
NOR2_X1 \myidu/_1160_ ( .A1(\myidu/_0163_ ), .A2(\myidu/_0164_ ), .ZN(\myidu/_0336_ ) );
NOR2_X1 \myidu/_1161_ ( .A1(\myidu/_0162_ ), .A2(\myidu/_0165_ ), .ZN(\myidu/_0337_ ) );
AND2_X1 \myidu/_1162_ ( .A1(\myidu/_0336_ ), .A2(\myidu/_0337_ ), .ZN(\myidu/_0338_ ) );
INV_X1 \myidu/_1163_ ( .A(\myidu/_0168_ ), .ZN(\myidu/_0339_ ) );
NOR2_X1 \myidu/_1164_ ( .A1(\myidu/_0169_ ), .A2(\myidu/_0170_ ), .ZN(\myidu/_0340_ ) );
AND4_X1 \myidu/_1165_ ( .A1(\myidu/_0167_ ), .A2(\myidu/_0338_ ), .A3(\myidu/_0339_ ), .A4(\myidu/_0340_ ), .ZN(\myidu/_0341_ ) );
NAND3_X1 \myidu/_1166_ ( .A1(\myidu/_0282_ ), .A2(\myidu/_0272_ ), .A3(\myidu/_0283_ ), .ZN(\myidu/_0342_ ) );
NOR2_X1 \myidu/_1167_ ( .A1(\myidu/_0342_ ), .A2(\myidu/_0171_ ), .ZN(\myidu/_0343_ ) );
NOR2_X1 \myidu/_1168_ ( .A1(\myidu/_0179_ ), .A2(\myidu/_0178_ ), .ZN(\myidu/_0344_ ) );
AND2_X1 \myidu/_1169_ ( .A1(\myidu/_0271_ ), .A2(\myidu/_0344_ ), .ZN(\myidu/_0345_ ) );
AND2_X1 \myidu/_1170_ ( .A1(\myidu/_0343_ ), .A2(\myidu/_0345_ ), .ZN(\myidu/_0346_ ) );
AND2_X1 \myidu/_1171_ ( .A1(\myidu/_0341_ ), .A2(\myidu/_0346_ ), .ZN(\myidu/_0347_ ) );
NOR2_X1 \myidu/_1172_ ( .A1(\myidu/_0192_ ), .A2(\myidu/_0184_ ), .ZN(\myidu/_0348_ ) );
NAND4_X1 \myidu/_1173_ ( .A1(\myidu/_0348_ ), .A2(\myidu/_0202_ ), .A3(\myidu/_0300_ ), .A4(\myidu/_0203_ ), .ZN(\myidu/_0349_ ) );
NOR2_X1 \myidu/_1174_ ( .A1(\myidu/_0186_ ), .A2(\myidu/_0156_ ), .ZN(\myidu/_0350_ ) );
INV_X1 \myidu/_1175_ ( .A(\myidu/_0185_ ), .ZN(\myidu/_0351_ ) );
INV_X1 \myidu/_1176_ ( .A(\myidu/_0157_ ), .ZN(\myidu/_0352_ ) );
NAND3_X1 \myidu/_1177_ ( .A1(\myidu/_0350_ ), .A2(\myidu/_0351_ ), .A3(\myidu/_0352_ ), .ZN(\myidu/_0353_ ) );
INV_X1 \myidu/_1178_ ( .A(\myidu/_0161_ ), .ZN(\myidu/_0354_ ) );
NAND4_X1 \myidu/_1179_ ( .A1(\myidu/_0354_ ), .A2(\myidu/_0200_ ), .A3(\myidu/_0226_ ), .A4(\myidu/_0208_ ), .ZN(\myidu/_0355_ ) );
NOR3_X1 \myidu/_1180_ ( .A1(\myidu/_0349_ ), .A2(\myidu/_0353_ ), .A3(\myidu/_0355_ ), .ZN(\myidu/_0356_ ) );
AND2_X1 \myidu/_1181_ ( .A1(\myidu/_0347_ ), .A2(\myidu/_0356_ ), .ZN(\myidu/_0357_ ) );
AND2_X1 \myidu/_1182_ ( .A1(\myidu/_0196_ ), .A2(\myidu/_0180_ ), .ZN(\myidu/_0358_ ) );
INV_X1 \myidu/_1183_ ( .A(\myidu/_0358_ ), .ZN(\myidu/_0359_ ) );
BUF_X2 \myidu/_1184_ ( .A(\myidu/_0194_ ), .Z(\myidu/_0360_ ) );
NAND4_X1 \myidu/_1185_ ( .A1(\myidu/_0360_ ), .A2(\myidu/_0215_ ), .A3(\myidu/_0192_ ), .A4(\myidu/_0158_ ), .ZN(\myidu/_0361_ ) );
NOR2_X1 \myidu/_1186_ ( .A1(\myidu/_0359_ ), .A2(\myidu/_0361_ ), .ZN(\myidu/_0362_ ) );
NOR2_X1 \myidu/_1187_ ( .A1(\myidu/_0357_ ), .A2(\myidu/_0362_ ), .ZN(\myidu/_0363_ ) );
INV_X1 \myidu/_1188_ ( .A(\myidu/_0194_ ), .ZN(\myidu/_0364_ ) );
NOR4_X1 \myidu/_1189_ ( .A1(\myidu/_0353_ ), .A2(\myidu/_0364_ ), .A3(\myidu/_0161_ ), .A4(\myidu/_0184_ ), .ZN(\myidu/_0365_ ) );
AND2_X1 \myidu/_1190_ ( .A1(\myidu/_0365_ ), .A2(\myidu/_0232_ ), .ZN(\myidu/_0366_ ) );
AND2_X1 \myidu/_1191_ ( .A1(\myidu/_0338_ ), .A2(\myidu/_0340_ ), .ZN(\myidu/_0367_ ) );
INV_X1 \myidu/_1192_ ( .A(\myidu/_0167_ ), .ZN(\myidu/_0368_ ) );
AND3_X1 \myidu/_1193_ ( .A1(\myidu/_0367_ ), .A2(\myidu/_0368_ ), .A3(\myidu/_0339_ ), .ZN(\myidu/_0369_ ) );
AND2_X1 \myidu/_1194_ ( .A1(\myidu/_0369_ ), .A2(\myidu/_0346_ ), .ZN(\myidu/_0370_ ) );
AND4_X1 \myidu/_1195_ ( .A1(\myidu/_0368_ ), .A2(\myidu/_0168_ ), .A3(\myidu/_0176_ ), .A4(\myidu/_0175_ ), .ZN(\myidu/_0371_ ) );
AND3_X1 \myidu/_1196_ ( .A1(\myidu/_0371_ ), .A2(\myidu/_0344_ ), .A3(\myidu/_0340_ ), .ZN(\myidu/_0372_ ) );
AND3_X1 \myidu/_1197_ ( .A1(\myidu/_0372_ ), .A2(\myidu/_0343_ ), .A3(\myidu/_0338_ ), .ZN(\myidu/_0373_ ) );
OAI21_X1 \myidu/_1198_ ( .A(\myidu/_0366_ ), .B1(\myidu/_0370_ ), .B2(\myidu/_0373_ ), .ZN(\myidu/_0374_ ) );
AND3_X1 \myidu/_1199_ ( .A1(\myidu/_0196_ ), .A2(\myidu/_0197_ ), .A3(\myidu/_0192_ ), .ZN(\myidu/_0375_ ) );
AND2_X1 \myidu/_1200_ ( .A1(\myidu/_0375_ ), .A2(\myidu/_0181_ ), .ZN(\myidu/_0376_ ) );
INV_X1 \myidu/_1201_ ( .A(\myidu/_0376_ ), .ZN(\myidu/_0377_ ) );
AND4_X4 \myidu/_1202_ ( .A1(\myidu/_0268_ ), .A2(\myidu/_0363_ ), .A3(\myidu/_0374_ ), .A4(\myidu/_0377_ ), .ZN(\myidu/_0378_ ) );
AND2_X1 \myidu/_1203_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0279_ ), .ZN(\myidu/_0379_ ) );
AOI22_X1 \myidu/_1204_ ( .A1(\myidu/_0379_ ), .A2(\myidu/_0299_ ), .B1(\myidu/_0280_ ), .B2(\myidu/_0293_ ), .ZN(\myidu/_0380_ ) );
AND4_X1 \myidu/_1205_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0279_ ), .A3(\myidu/_0269_ ), .A4(\myidu/_0298_ ), .ZN(\myidu/_0381_ ) );
AOI21_X1 \myidu/_1206_ ( .A(\myidu/_0381_ ), .B1(\myidu/_0379_ ), .B2(\myidu/_0305_ ), .ZN(\myidu/_0382_ ) );
NAND3_X1 \myidu/_1207_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0293_ ), .A3(\myidu/_0279_ ), .ZN(\myidu/_0383_ ) );
NAND3_X1 \myidu/_1208_ ( .A1(\myidu/_0285_ ), .A2(\myidu/_0204_ ), .A3(\myidu/_0279_ ), .ZN(\myidu/_0384_ ) );
AND2_X1 \myidu/_1209_ ( .A1(\myidu/_0383_ ), .A2(\myidu/_0384_ ), .ZN(\myidu/_0385_ ) );
NAND3_X1 \myidu/_1210_ ( .A1(\myidu/_0380_ ), .A2(\myidu/_0382_ ), .A3(\myidu/_0385_ ), .ZN(\myidu/_0386_ ) );
NAND3_X1 \myidu/_1211_ ( .A1(\myidu/_0281_ ), .A2(\myidu/_0286_ ), .A3(\myidu/_0288_ ), .ZN(\myidu/_0387_ ) );
NOR3_X4 \myidu/_1212_ ( .A1(\myidu/_0386_ ), .A2(\myidu/_0387_ ), .A3(\myidu/_0332_ ), .ZN(\myidu/_0388_ ) );
AND2_X1 \myidu/_1213_ ( .A1(\myidu/_0378_ ), .A2(\myidu/_0388_ ), .ZN(\myidu/_0389_ ) );
AND3_X1 \myidu/_1214_ ( .A1(\myidu/_0205_ ), .A2(\myidu/_0182_ ), .A3(\myidu/_0183_ ), .ZN(\myidu/_0390_ ) );
AND2_X1 \myidu/_1215_ ( .A1(\myidu/_0358_ ), .A2(\myidu/_0390_ ), .ZN(\myidu/_0391_ ) );
INV_X1 \myidu/_1216_ ( .A(\myidu/_0391_ ), .ZN(\myidu/_0392_ ) );
AOI21_X1 \myidu/_1217_ ( .A(\myidu/_0335_ ), .B1(\myidu/_0389_ ), .B2(\myidu/_0392_ ), .ZN(\myidu/_0393_ ) );
OAI21_X1 \myidu/_1218_ ( .A(\myidu/_0334_ ), .B1(\myidu/_0393_ ), .B2(\myidu/_0368_ ), .ZN(\myidu/_0394_ ) );
NAND3_X1 \myidu/_1219_ ( .A1(\myidu/_0224_ ), .A2(\myidu/_0229_ ), .A3(\myidu/_0392_ ), .ZN(\myidu/_0395_ ) );
NAND2_X4 \myidu/_1220_ ( .A1(\myidu/_0378_ ), .A2(\myidu/_0388_ ), .ZN(\myidu/_0396_ ) );
INV_X1 \myidu/_1221_ ( .A(\myidu/_0295_ ), .ZN(\myidu/_0397_ ) );
NOR3_X4 \myidu/_1222_ ( .A1(\myidu/_0395_ ), .A2(\myidu/_0396_ ), .A3(\myidu/_0397_ ), .ZN(\myidu/_0398_ ) );
INV_X1 \myidu/_1223_ ( .A(\myidu/_0319_ ), .ZN(\myidu/_0399_ ) );
NOR2_X4 \myidu/_1224_ ( .A1(\myidu/_0398_ ), .A2(\myidu/_0399_ ), .ZN(\myidu/_0400_ ) );
AND2_X4 \myidu/_1225_ ( .A1(\myidu/_0400_ ), .A2(\myidu/_0322_ ), .ZN(\myidu/_0401_ ) );
BUF_X8 \myidu/_1226_ ( .A(\myidu/_0401_ ), .Z(\myidu/_0402_ ) );
MUX2_X1 \myidu/_1227_ ( .A(\myidu/_0123_ ), .B(\myidu/_0394_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0008_ ) );
AND2_X1 \myidu/_1228_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0162_ ), .ZN(\myidu/_0403_ ) );
INV_X1 \myidu/_1229_ ( .A(\myidu/_0268_ ), .ZN(\myidu/_0404_ ) );
AOI21_X1 \myidu/_1230_ ( .A(\myidu/_0403_ ), .B1(\myidu/_0404_ ), .B2(\myidu/_0185_ ), .ZN(\myidu/_0405_ ) );
OAI21_X1 \myidu/_1231_ ( .A(\myidu/_0405_ ), .B1(\myidu/_0396_ ), .B2(\myidu/_0339_ ), .ZN(\myidu/_0406_ ) );
MUX2_X1 \myidu/_1232_ ( .A(\myidu/_0134_ ), .B(\myidu/_0406_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0009_ ) );
AND2_X1 \myidu/_1233_ ( .A1(\myidu/_0332_ ), .A2(\myidu/_0163_ ), .ZN(\myidu/_0407_ ) );
AOI21_X1 \myidu/_1234_ ( .A(\myidu/_0407_ ), .B1(\myidu/_0404_ ), .B2(\myidu/_0186_ ), .ZN(\myidu/_0408_ ) );
INV_X1 \myidu/_1235_ ( .A(\myidu/_0169_ ), .ZN(\myidu/_0409_ ) );
OAI21_X1 \myidu/_1236_ ( .A(\myidu/_0408_ ), .B1(\myidu/_0396_ ), .B2(\myidu/_0409_ ), .ZN(\myidu/_0410_ ) );
MUX2_X1 \myidu/_1237_ ( .A(\myidu/_0145_ ), .B(\myidu/_0410_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0010_ ) );
AND2_X1 \myidu/_1238_ ( .A1(\myidu/_0332_ ), .A2(\myidu/_0164_ ), .ZN(\myidu/_0411_ ) );
AOI21_X1 \myidu/_1239_ ( .A(\myidu/_0411_ ), .B1(\myidu/_0404_ ), .B2(\myidu/_0156_ ), .ZN(\myidu/_0412_ ) );
INV_X1 \myidu/_1240_ ( .A(\myidu/_0170_ ), .ZN(\myidu/_0413_ ) );
OAI21_X1 \myidu/_1241_ ( .A(\myidu/_0412_ ), .B1(\myidu/_0396_ ), .B2(\myidu/_0413_ ), .ZN(\myidu/_0414_ ) );
MUX2_X1 \myidu/_1242_ ( .A(\myidu/_0148_ ), .B(\myidu/_0414_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0011_ ) );
AND2_X1 \myidu/_1243_ ( .A1(\myidu/_0332_ ), .A2(\myidu/_0165_ ), .ZN(\myidu/_0415_ ) );
AOI21_X1 \myidu/_1244_ ( .A(\myidu/_0415_ ), .B1(\myidu/_0404_ ), .B2(\myidu/_0157_ ), .ZN(\myidu/_0416_ ) );
INV_X1 \myidu/_1245_ ( .A(\myidu/_0171_ ), .ZN(\myidu/_0417_ ) );
OAI21_X1 \myidu/_1246_ ( .A(\myidu/_0416_ ), .B1(\myidu/_0396_ ), .B2(\myidu/_0417_ ), .ZN(\myidu/_0418_ ) );
MUX2_X1 \myidu/_1247_ ( .A(\myidu/_0149_ ), .B(\myidu/_0418_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0012_ ) );
OR2_X1 \myidu/_1248_ ( .A1(\myidu/_0395_ ), .A2(\myidu/_0404_ ), .ZN(\myidu/_0419_ ) );
AND2_X1 \myidu/_1249_ ( .A1(\myidu/_0419_ ), .A2(\myidu/_0172_ ), .ZN(\myidu/_0420_ ) );
MUX2_X1 \myidu/_1250_ ( .A(\myidu/_0150_ ), .B(\myidu/_0420_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0013_ ) );
AND2_X1 \myidu/_1251_ ( .A1(\myidu/_0419_ ), .A2(\myidu/_0173_ ), .ZN(\myidu/_0421_ ) );
MUX2_X1 \myidu/_1252_ ( .A(\myidu/_0151_ ), .B(\myidu/_0421_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0014_ ) );
AND2_X1 \myidu/_1253_ ( .A1(\myidu/_0419_ ), .A2(\myidu/_0174_ ), .ZN(\myidu/_0422_ ) );
MUX2_X1 \myidu/_1254_ ( .A(\myidu/_0152_ ), .B(\myidu/_0422_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0015_ ) );
AND2_X1 \myidu/_1255_ ( .A1(\myidu/_0419_ ), .A2(\myidu/_0175_ ), .ZN(\myidu/_0423_ ) );
MUX2_X1 \myidu/_1256_ ( .A(\myidu/_0153_ ), .B(\myidu/_0423_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0016_ ) );
AND2_X1 \myidu/_1257_ ( .A1(\myidu/_0419_ ), .A2(\myidu/_0176_ ), .ZN(\myidu/_0424_ ) );
MUX2_X1 \myidu/_1258_ ( .A(\myidu/_0154_ ), .B(\myidu/_0424_ ), .S(\myidu/_0402_ ), .Z(\myidu/_0017_ ) );
AND2_X1 \myidu/_1259_ ( .A1(\myidu/_0419_ ), .A2(\myidu/_0178_ ), .ZN(\myidu/_0425_ ) );
BUF_X8 \myidu/_1260_ ( .A(\myidu/_0401_ ), .Z(\myidu/_0426_ ) );
MUX2_X1 \myidu/_1261_ ( .A(\myidu/_0124_ ), .B(\myidu/_0425_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0018_ ) );
AOI21_X1 \myidu/_1262_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0261_ ), .B2(\myidu/_0262_ ), .ZN(\myidu/_0427_ ) );
AOI221_X4 \myidu/_1263_ ( .A(\myidu/_0427_ ), .B1(\myidu/_0167_ ), .B2(\myidu/_0391_ ), .C1(\myidu/_0184_ ), .C2(\myidu/_0267_ ), .ZN(\myidu/_0428_ ) );
BUF_X4 \myidu/_1264_ ( .A(\myidu/_0290_ ), .Z(\myidu/_0429_ ) );
OAI21_X1 \myidu/_1265_ ( .A(\myidu/_0428_ ), .B1(\myidu/_0230_ ), .B2(\myidu/_0429_ ), .ZN(\myidu/_0430_ ) );
MUX2_X1 \myidu/_1266_ ( .A(\myidu/_0125_ ), .B(\myidu/_0430_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0019_ ) );
AOI21_X1 \myidu/_1267_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0224_ ), .B2(\myidu/_0229_ ), .ZN(\myidu/_0431_ ) );
NOR2_X1 \myidu/_1268_ ( .A1(\myidu/_0268_ ), .A2(\myidu/_0290_ ), .ZN(\myidu/_0432_ ) );
NOR2_X1 \myidu/_1269_ ( .A1(\myidu/_0431_ ), .A2(\myidu/_0432_ ), .ZN(\myidu/_0433_ ) );
NOR2_X2 \myidu/_1270_ ( .A1(\myidu/_0376_ ), .A2(\myidu/_0391_ ), .ZN(\myidu/_0434_ ) );
OAI21_X1 \myidu/_1271_ ( .A(\myidu/_0433_ ), .B1(\myidu/_0200_ ), .B2(\myidu/_0434_ ), .ZN(\myidu/_0435_ ) );
MUX2_X1 \myidu/_1272_ ( .A(\myidu/_0126_ ), .B(\myidu/_0435_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0020_ ) );
OAI21_X1 \myidu/_1273_ ( .A(\myidu/_0433_ ), .B1(\myidu/_0208_ ), .B2(\myidu/_0434_ ), .ZN(\myidu/_0436_ ) );
MUX2_X1 \myidu/_1274_ ( .A(\myidu/_0127_ ), .B(\myidu/_0436_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0021_ ) );
OAI21_X1 \myidu/_1275_ ( .A(\myidu/_0433_ ), .B1(\myidu/_0226_ ), .B2(\myidu/_0434_ ), .ZN(\myidu/_0437_ ) );
MUX2_X1 \myidu/_1276_ ( .A(\myidu/_0128_ ), .B(\myidu/_0437_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0022_ ) );
OAI21_X1 \myidu/_1277_ ( .A(\myidu/_0433_ ), .B1(\myidu/_0354_ ), .B2(\myidu/_0434_ ), .ZN(\myidu/_0438_ ) );
MUX2_X1 \myidu/_1278_ ( .A(\myidu/_0129_ ), .B(\myidu/_0438_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0023_ ) );
CLKBUF_X2 \myidu/_1279_ ( .A(\myidu/_0432_ ), .Z(\myidu/_0439_ ) );
INV_X1 \myidu/_1280_ ( .A(\myidu/_0434_ ), .ZN(\myidu/_0440_ ) );
AND2_X1 \myidu/_1281_ ( .A1(\myidu/_0440_ ), .A2(\myidu/_0162_ ), .ZN(\myidu/_0441_ ) );
OR3_X1 \myidu/_1282_ ( .A1(\myidu/_0431_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0441_ ), .ZN(\myidu/_0442_ ) );
MUX2_X1 \myidu/_1283_ ( .A(\myidu/_0130_ ), .B(\myidu/_0442_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0024_ ) );
AND2_X1 \myidu/_1284_ ( .A1(\myidu/_0440_ ), .A2(\myidu/_0163_ ), .ZN(\myidu/_0443_ ) );
OR3_X1 \myidu/_1285_ ( .A1(\myidu/_0431_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0443_ ), .ZN(\myidu/_0444_ ) );
MUX2_X1 \myidu/_1286_ ( .A(\myidu/_0131_ ), .B(\myidu/_0444_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0025_ ) );
AND2_X1 \myidu/_1287_ ( .A1(\myidu/_0440_ ), .A2(\myidu/_0164_ ), .ZN(\myidu/_0445_ ) );
OR3_X1 \myidu/_1288_ ( .A1(\myidu/_0431_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0445_ ), .ZN(\myidu/_0446_ ) );
MUX2_X1 \myidu/_1289_ ( .A(\myidu/_0132_ ), .B(\myidu/_0446_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0026_ ) );
AND2_X1 \myidu/_1290_ ( .A1(\myidu/_0440_ ), .A2(\myidu/_0165_ ), .ZN(\myidu/_0447_ ) );
OR3_X1 \myidu/_1291_ ( .A1(\myidu/_0431_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0447_ ), .ZN(\myidu/_0448_ ) );
MUX2_X1 \myidu/_1292_ ( .A(\myidu/_0133_ ), .B(\myidu/_0448_ ), .S(\myidu/_0426_ ), .Z(\myidu/_0027_ ) );
AND2_X2 \myidu/_1293_ ( .A1(\myidu/_0395_ ), .A2(\myidu/_0179_ ), .ZN(\myidu/_0449_ ) );
CLKBUF_X2 \myidu/_1294_ ( .A(\myidu/_0449_ ), .Z(\myidu/_0450_ ) );
CLKBUF_X2 \myidu/_1295_ ( .A(\myidu/_0375_ ), .Z(\myidu/_0451_ ) );
AND3_X1 \myidu/_1296_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0167_ ), .A3(\myidu/_0181_ ), .ZN(\myidu/_0452_ ) );
OR3_X1 \myidu/_1297_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0452_ ), .ZN(\myidu/_0453_ ) );
BUF_X8 \myidu/_1298_ ( .A(\myidu/_0401_ ), .Z(\myidu/_0454_ ) );
MUX2_X1 \myidu/_1299_ ( .A(\myidu/_0135_ ), .B(\myidu/_0453_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0028_ ) );
AND3_X1 \myidu/_1300_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0168_ ), .A3(\myidu/_0181_ ), .ZN(\myidu/_0455_ ) );
OR3_X1 \myidu/_1301_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0455_ ), .ZN(\myidu/_0456_ ) );
MUX2_X1 \myidu/_1302_ ( .A(\myidu/_0136_ ), .B(\myidu/_0456_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0029_ ) );
AND3_X1 \myidu/_1303_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0169_ ), .A3(\myidu/_0181_ ), .ZN(\myidu/_0457_ ) );
OR3_X1 \myidu/_1304_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0457_ ), .ZN(\myidu/_0458_ ) );
MUX2_X1 \myidu/_1305_ ( .A(\myidu/_0137_ ), .B(\myidu/_0458_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0030_ ) );
AND3_X1 \myidu/_1306_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0170_ ), .A3(\myidu/_0181_ ), .ZN(\myidu/_0459_ ) );
OR3_X1 \myidu/_1307_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0459_ ), .ZN(\myidu/_0460_ ) );
MUX2_X1 \myidu/_1308_ ( .A(\myidu/_0138_ ), .B(\myidu/_0460_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0031_ ) );
AND3_X1 \myidu/_1309_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0171_ ), .A3(\myidu/_0181_ ), .ZN(\myidu/_0461_ ) );
OR3_X1 \myidu/_1310_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0461_ ), .ZN(\myidu/_0462_ ) );
MUX2_X1 \myidu/_1311_ ( .A(\myidu/_0139_ ), .B(\myidu/_0462_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0032_ ) );
AND3_X1 \myidu/_1312_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0172_ ), .ZN(\myidu/_0463_ ) );
OR3_X1 \myidu/_1313_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0439_ ), .A3(\myidu/_0463_ ), .ZN(\myidu/_0464_ ) );
MUX2_X1 \myidu/_1314_ ( .A(\myidu/_0140_ ), .B(\myidu/_0464_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0033_ ) );
AND3_X1 \myidu/_1315_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0173_ ), .ZN(\myidu/_0465_ ) );
OR3_X1 \myidu/_1316_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0432_ ), .A3(\myidu/_0465_ ), .ZN(\myidu/_0466_ ) );
MUX2_X1 \myidu/_1317_ ( .A(\myidu/_0141_ ), .B(\myidu/_0466_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0034_ ) );
AND3_X1 \myidu/_1318_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0174_ ), .ZN(\myidu/_0467_ ) );
OR3_X1 \myidu/_1319_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0432_ ), .A3(\myidu/_0467_ ), .ZN(\myidu/_0468_ ) );
MUX2_X1 \myidu/_1320_ ( .A(\myidu/_0142_ ), .B(\myidu/_0468_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0035_ ) );
AND3_X1 \myidu/_1321_ ( .A1(\myidu/_0451_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0175_ ), .ZN(\myidu/_0469_ ) );
OR3_X1 \myidu/_1322_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0432_ ), .A3(\myidu/_0469_ ), .ZN(\myidu/_0470_ ) );
MUX2_X1 \myidu/_1323_ ( .A(\myidu/_0143_ ), .B(\myidu/_0470_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0036_ ) );
AND3_X1 \myidu/_1324_ ( .A1(\myidu/_0375_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0176_ ), .ZN(\myidu/_0471_ ) );
OR3_X1 \myidu/_1325_ ( .A1(\myidu/_0449_ ), .A2(\myidu/_0432_ ), .A3(\myidu/_0471_ ), .ZN(\myidu/_0472_ ) );
MUX2_X1 \myidu/_1326_ ( .A(\myidu/_0144_ ), .B(\myidu/_0472_ ), .S(\myidu/_0454_ ), .Z(\myidu/_0037_ ) );
AND3_X1 \myidu/_1327_ ( .A1(\myidu/_0375_ ), .A2(\myidu/_0181_ ), .A3(\myidu/_0178_ ), .ZN(\myidu/_0473_ ) );
OR3_X1 \myidu/_1328_ ( .A1(\myidu/_0449_ ), .A2(\myidu/_0432_ ), .A3(\myidu/_0473_ ), .ZN(\myidu/_0474_ ) );
MUX2_X1 \myidu/_1329_ ( .A(\myidu/_0146_ ), .B(\myidu/_0474_ ), .S(\myidu/_0401_ ), .Z(\myidu/_0038_ ) );
AOI21_X1 \myidu/_1330_ ( .A(\myidu/_0429_ ), .B1(\myidu/_0268_ ), .B2(\myidu/_0377_ ), .ZN(\myidu/_0475_ ) );
OR2_X1 \myidu/_1331_ ( .A1(\myidu/_0450_ ), .A2(\myidu/_0475_ ), .ZN(\myidu/_0476_ ) );
MUX2_X1 \myidu/_1332_ ( .A(\myidu/_0147_ ), .B(\myidu/_0476_ ), .S(\myidu/_0401_ ), .Z(\myidu/_0039_ ) );
AND2_X2 \myidu/_1333_ ( .A1(\myidu/_0319_ ), .A2(\myidu/_0322_ ), .ZN(\myidu/_0477_ ) );
BUF_X4 \myidu/_1334_ ( .A(\myidu/_0477_ ), .Z(\myidu/_0478_ ) );
MUX2_X1 \myidu/_1335_ ( .A(\myidu/_0740_ ), .B(\myidu/_0708_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0049_ ) );
MUX2_X1 \myidu/_1336_ ( .A(\myidu/_0751_ ), .B(\myidu/_0719_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0050_ ) );
MUX2_X1 \myidu/_1337_ ( .A(\myidu/_0762_ ), .B(\myidu/_0730_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0051_ ) );
MUX2_X1 \myidu/_1338_ ( .A(\myidu/_0765_ ), .B(\myidu/_0733_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0052_ ) );
MUX2_X1 \myidu/_1339_ ( .A(\myidu/_0766_ ), .B(\myidu/_0734_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0053_ ) );
MUX2_X1 \myidu/_1340_ ( .A(\myidu/_0767_ ), .B(\myidu/_0735_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0054_ ) );
MUX2_X1 \myidu/_1341_ ( .A(\myidu/_0768_ ), .B(\myidu/_0736_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0055_ ) );
MUX2_X1 \myidu/_1342_ ( .A(\myidu/_0769_ ), .B(\myidu/_0737_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0056_ ) );
MUX2_X1 \myidu/_1343_ ( .A(\myidu/_0770_ ), .B(\myidu/_0738_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0057_ ) );
MUX2_X1 \myidu/_1344_ ( .A(\myidu/_0771_ ), .B(\myidu/_0739_ ), .S(\myidu/_0478_ ), .Z(\myidu/_0058_ ) );
BUF_X4 \myidu/_1345_ ( .A(\myidu/_0477_ ), .Z(\myidu/_0479_ ) );
MUX2_X1 \myidu/_1346_ ( .A(\myidu/_0741_ ), .B(\myidu/_0709_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0059_ ) );
MUX2_X1 \myidu/_1347_ ( .A(\myidu/_0742_ ), .B(\myidu/_0710_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0060_ ) );
MUX2_X1 \myidu/_1348_ ( .A(\myidu/_0743_ ), .B(\myidu/_0711_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0061_ ) );
MUX2_X1 \myidu/_1349_ ( .A(\myidu/_0744_ ), .B(\myidu/_0712_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0062_ ) );
MUX2_X1 \myidu/_1350_ ( .A(\myidu/_0745_ ), .B(\myidu/_0713_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0063_ ) );
MUX2_X1 \myidu/_1351_ ( .A(\myidu/_0746_ ), .B(\myidu/_0714_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0064_ ) );
MUX2_X1 \myidu/_1352_ ( .A(\myidu/_0747_ ), .B(\myidu/_0715_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0065_ ) );
MUX2_X1 \myidu/_1353_ ( .A(\myidu/_0748_ ), .B(\myidu/_0716_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0066_ ) );
MUX2_X1 \myidu/_1354_ ( .A(\myidu/_0749_ ), .B(\myidu/_0717_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0067_ ) );
MUX2_X1 \myidu/_1355_ ( .A(\myidu/_0750_ ), .B(\myidu/_0718_ ), .S(\myidu/_0479_ ), .Z(\myidu/_0068_ ) );
BUF_X4 \myidu/_1356_ ( .A(\myidu/_0477_ ), .Z(\myidu/_0480_ ) );
MUX2_X1 \myidu/_1357_ ( .A(\myidu/_0752_ ), .B(\myidu/_0720_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0069_ ) );
MUX2_X1 \myidu/_1358_ ( .A(\myidu/_0753_ ), .B(\myidu/_0721_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0070_ ) );
MUX2_X1 \myidu/_1359_ ( .A(\myidu/_0754_ ), .B(\myidu/_0722_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0071_ ) );
MUX2_X1 \myidu/_1360_ ( .A(\myidu/_0755_ ), .B(\myidu/_0723_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0072_ ) );
MUX2_X1 \myidu/_1361_ ( .A(\myidu/_0756_ ), .B(\myidu/_0724_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0073_ ) );
MUX2_X1 \myidu/_1362_ ( .A(\myidu/_0757_ ), .B(\myidu/_0725_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0074_ ) );
MUX2_X1 \myidu/_1363_ ( .A(\myidu/_0758_ ), .B(\myidu/_0726_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0075_ ) );
MUX2_X1 \myidu/_1364_ ( .A(\myidu/_0759_ ), .B(\myidu/_0727_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0076_ ) );
MUX2_X1 \myidu/_1365_ ( .A(\myidu/_0760_ ), .B(\myidu/_0728_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0077_ ) );
MUX2_X1 \myidu/_1366_ ( .A(\myidu/_0761_ ), .B(\myidu/_0729_ ), .S(\myidu/_0480_ ), .Z(\myidu/_0078_ ) );
MUX2_X1 \myidu/_1367_ ( .A(\myidu/_0763_ ), .B(\myidu/_0731_ ), .S(\myidu/_0477_ ), .Z(\myidu/_0079_ ) );
MUX2_X1 \myidu/_1368_ ( .A(\myidu/_0764_ ), .B(\myidu/_0732_ ), .S(\myidu/_0477_ ), .Z(\myidu/_0080_ ) );
NOR2_X1 \myidu/_1369_ ( .A1(\myidu/_0326_ ), .A2(\myidu/_0801_ ), .ZN(\myidu/_0481_ ) );
OAI221_X1 \myidu/_1370_ ( .A(\myidu/_0323_ ), .B1(\myidu/_0320_ ), .B2(\myidu/_0790_ ), .C1(\myidu/_0481_ ), .C2(\myidu/_0188_ ), .ZN(\myidu/_0482_ ) );
INV_X1 \myidu/_1371_ ( .A(\myidu/_0362_ ), .ZN(\myidu/_0483_ ) );
BUF_X4 \myidu/_1372_ ( .A(\myidu/_0320_ ), .Z(\myidu/_0484_ ) );
AOI21_X1 \myidu/_1373_ ( .A(\myidu/_0482_ ), .B1(\myidu/_0483_ ), .B2(\myidu/_0484_ ), .ZN(\myidu/_0040_ ) );
BUF_X2 \myidu/_1374_ ( .A(\myidu/_0211_ ), .Z(\myidu/_0485_ ) );
CLKBUF_X2 \myidu/_1375_ ( .A(\myidu/_0485_ ), .Z(\myidu/_0486_ ) );
AND3_X1 \myidu/_1376_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0221_ ), .A3(\myidu/_0234_ ), .ZN(\myidu/_0487_ ) );
OR2_X1 \myidu/_1377_ ( .A1(\myidu/_0357_ ), .A2(\myidu/_0487_ ), .ZN(\myidu/_0488_ ) );
NOR2_X1 \myidu/_1378_ ( .A1(\myidu/_0226_ ), .A2(\myidu/_0159_ ), .ZN(\myidu/_0489_ ) );
AOI221_X4 \myidu/_1379_ ( .A(\myidu/_0488_ ), .B1(\myidu/_0489_ ), .B2(\myidu/_0235_ ), .C1(\myidu/_0221_ ), .C2(\myidu/_0232_ ), .ZN(\myidu/_0490_ ) );
NAND4_X1 \myidu/_1380_ ( .A1(\myidu/_0191_ ), .A2(\myidu/_0196_ ), .A3(\myidu/_0193_ ), .A4(\myidu/_0197_ ), .ZN(\myidu/_0491_ ) );
NOR2_X1 \myidu/_1381_ ( .A1(\myidu/_0491_ ), .A2(\myidu/_0364_ ), .ZN(\myidu/_0492_ ) );
INV_X1 \myidu/_1382_ ( .A(\myidu/_0492_ ), .ZN(\myidu/_0493_ ) );
AND3_X1 \myidu/_1383_ ( .A1(\myidu/_0297_ ), .A2(\myidu/_0303_ ), .A3(\myidu/_0191_ ), .ZN(\myidu/_0494_ ) );
NAND2_X1 \myidu/_1384_ ( .A1(\myidu/_0494_ ), .A2(\myidu/_0209_ ), .ZN(\myidu/_0495_ ) );
AND2_X1 \myidu/_1385_ ( .A1(\myidu/_0494_ ), .A2(\myidu/_0360_ ), .ZN(\myidu/_0496_ ) );
NAND4_X1 \myidu/_1386_ ( .A1(\myidu/_0308_ ), .A2(\myidu/_0191_ ), .A3(\myidu/_0202_ ), .A4(\myidu/_0203_ ), .ZN(\myidu/_0497_ ) );
NOR2_X1 \myidu/_1387_ ( .A1(\myidu/_0497_ ), .A2(\myidu/_0364_ ), .ZN(\myidu/_0498_ ) );
OR2_X1 \myidu/_1388_ ( .A1(\myidu/_0496_ ), .A2(\myidu/_0498_ ), .ZN(\myidu/_0499_ ) );
AND4_X1 \myidu/_1389_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0275_ ), .A3(\myidu/_0287_ ), .A4(\myidu/_0206_ ), .ZN(\myidu/_0500_ ) );
INV_X1 \myidu/_1390_ ( .A(\myidu/_0500_ ), .ZN(\myidu/_0501_ ) );
AND4_X1 \myidu/_1391_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0270_ ), .A3(\myidu/_0273_ ), .A4(\myidu/_0206_ ), .ZN(\myidu/_0502_ ) );
INV_X1 \myidu/_1392_ ( .A(\myidu/_0502_ ), .ZN(\myidu/_0503_ ) );
AOI21_X1 \myidu/_1393_ ( .A(\myidu/_0179_ ), .B1(\myidu/_0501_ ), .B2(\myidu/_0503_ ), .ZN(\myidu/_0504_ ) );
NOR2_X1 \myidu/_1394_ ( .A1(\myidu/_0499_ ), .A2(\myidu/_0504_ ), .ZN(\myidu/_0505_ ) );
AND3_X2 \myidu/_1395_ ( .A1(\myidu/_0485_ ), .A2(\myidu/_0303_ ), .A3(\myidu/_0215_ ), .ZN(\myidu/_0506_ ) );
NAND2_X1 \myidu/_1396_ ( .A1(\myidu/_0506_ ), .A2(\myidu/_0489_ ), .ZN(\myidu/_0507_ ) );
AND3_X1 \myidu/_1397_ ( .A1(\myidu/_0485_ ), .A2(\myidu/_0308_ ), .A3(\myidu/_0215_ ), .ZN(\myidu/_0508_ ) );
AND2_X1 \myidu/_1398_ ( .A1(\myidu/_0183_ ), .A2(\myidu/_0158_ ), .ZN(\myidu/_0509_ ) );
AND3_X1 \myidu/_1399_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0191_ ), .A3(\myidu/_0509_ ), .ZN(\myidu/_0510_ ) );
AOI22_X1 \myidu/_1400_ ( .A1(\myidu/_0489_ ), .A2(\myidu/_0508_ ), .B1(\myidu/_0510_ ), .B2(\myidu/_0360_ ), .ZN(\myidu/_0511_ ) );
AND4_X1 \myidu/_1401_ ( .A1(\myidu/_0495_ ), .A2(\myidu/_0505_ ), .A3(\myidu/_0507_ ), .A4(\myidu/_0511_ ), .ZN(\myidu/_0512_ ) );
AND3_X1 \myidu/_1402_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0191_ ), .A3(\myidu/_0193_ ), .ZN(\myidu/_0513_ ) );
OAI21_X1 \myidu/_1403_ ( .A(\myidu/_0221_ ), .B1(\myidu/_0513_ ), .B2(\myidu/_0510_ ), .ZN(\myidu/_0514_ ) );
NAND4_X1 \myidu/_1404_ ( .A1(\myidu/_0490_ ), .A2(\myidu/_0493_ ), .A3(\myidu/_0512_ ), .A4(\myidu/_0514_ ), .ZN(\myidu/_0515_ ) );
OAI21_X1 \myidu/_1405_ ( .A(\myidu/_0429_ ), .B1(\myidu/_0306_ ), .B2(\myidu/_0312_ ), .ZN(\myidu/_0516_ ) );
AND2_X1 \myidu/_1406_ ( .A1(\myidu/_0270_ ), .A2(\myidu/_0273_ ), .ZN(\myidu/_0517_ ) );
AND4_X1 \myidu/_1407_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0517_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0302_ ), .ZN(\myidu/_0518_ ) );
AND4_X1 \myidu/_1408_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0285_ ), .A3(\myidu/_0302_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0519_ ) );
OAI21_X1 \myidu/_1409_ ( .A(\myidu/_0429_ ), .B1(\myidu/_0518_ ), .B2(\myidu/_0519_ ), .ZN(\myidu/_0520_ ) );
NAND2_X1 \myidu/_1410_ ( .A1(\myidu/_0309_ ), .A2(\myidu/_0429_ ), .ZN(\myidu/_0521_ ) );
AND4_X1 \myidu/_1411_ ( .A1(\myidu/_0190_ ), .A2(\myidu/_0192_ ), .A3(\myidu/_0200_ ), .A4(\myidu/_0181_ ), .ZN(\myidu/_0522_ ) );
AND2_X2 \myidu/_1412_ ( .A1(\myidu/_0485_ ), .A2(\myidu/_0522_ ), .ZN(\myidu/_0523_ ) );
AOI22_X1 \myidu/_1413_ ( .A1(\myidu/_0207_ ), .A2(\myidu/_0221_ ), .B1(\myidu/_0489_ ), .B2(\myidu/_0523_ ), .ZN(\myidu/_0524_ ) );
NAND4_X1 \myidu/_1414_ ( .A1(\myidu/_0516_ ), .A2(\myidu/_0520_ ), .A3(\myidu/_0521_ ), .A4(\myidu/_0524_ ), .ZN(\myidu/_0525_ ) );
OAI21_X1 \myidu/_1415_ ( .A(\myidu/_0484_ ), .B1(\myidu/_0515_ ), .B2(\myidu/_0525_ ), .ZN(\myidu/_0526_ ) );
BUF_X4 \myidu/_1416_ ( .A(\myidu/_0399_ ), .Z(\myidu/_0527_ ) );
BUF_X4 \myidu/_1417_ ( .A(\myidu/_0527_ ), .Z(\myidu/_0528_ ) );
NAND2_X1 \myidu/_1418_ ( .A1(\myidu/_0528_ ), .A2(\myidu/_0793_ ), .ZN(\myidu/_0529_ ) );
AOI21_X1 \myidu/_1419_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0526_ ), .B2(\myidu/_0529_ ), .ZN(\myidu/_0041_ ) );
AND4_X1 \myidu/_1420_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0305_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0302_ ), .ZN(\myidu/_0530_ ) );
OAI21_X1 \myidu/_1421_ ( .A(\myidu/_0429_ ), .B1(\myidu/_0530_ ), .B2(\myidu/_0306_ ), .ZN(\myidu/_0531_ ) );
NAND2_X1 \myidu/_1422_ ( .A1(\myidu/_0518_ ), .A2(\myidu/_0429_ ), .ZN(\myidu/_0532_ ) );
NAND2_X1 \myidu/_1423_ ( .A1(\myidu/_0304_ ), .A2(\myidu/_0429_ ), .ZN(\myidu/_0533_ ) );
OAI21_X1 \myidu/_1424_ ( .A(\myidu/_0523_ ), .B1(\myidu/_0489_ ), .B2(\myidu/_0221_ ), .ZN(\myidu/_0534_ ) );
NAND4_X1 \myidu/_1425_ ( .A1(\myidu/_0531_ ), .A2(\myidu/_0532_ ), .A3(\myidu/_0533_ ), .A4(\myidu/_0534_ ), .ZN(\myidu/_0535_ ) );
NAND2_X1 \myidu/_1426_ ( .A1(\myidu/_0508_ ), .A2(\myidu/_0489_ ), .ZN(\myidu/_0536_ ) );
NAND3_X1 \myidu/_1427_ ( .A1(\myidu/_0216_ ), .A2(\myidu/_0486_ ), .A3(\myidu/_0360_ ), .ZN(\myidu/_0537_ ) );
AND3_X1 \myidu/_1428_ ( .A1(\myidu/_0495_ ), .A2(\myidu/_0536_ ), .A3(\myidu/_0537_ ), .ZN(\myidu/_0538_ ) );
AND4_X1 \myidu/_1429_ ( .A1(\myidu/_0204_ ), .A2(\myidu/_0275_ ), .A3(\myidu/_0270_ ), .A4(\myidu/_0206_ ), .ZN(\myidu/_0539_ ) );
OAI21_X1 \myidu/_1430_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0539_ ), .B2(\myidu/_0502_ ), .ZN(\myidu/_0540_ ) );
AOI22_X1 \myidu/_1431_ ( .A1(\myidu/_0513_ ), .A2(\myidu/_0160_ ), .B1(\myidu/_0232_ ), .B2(\myidu/_0159_ ), .ZN(\myidu/_0541_ ) );
AOI21_X1 \myidu/_1432_ ( .A(\myidu/_0498_ ), .B1(\myidu/_0302_ ), .B2(\myidu/_0451_ ), .ZN(\myidu/_0542_ ) );
NAND4_X1 \myidu/_1433_ ( .A1(\myidu/_0538_ ), .A2(\myidu/_0540_ ), .A3(\myidu/_0541_ ), .A4(\myidu/_0542_ ), .ZN(\myidu/_0543_ ) );
OAI21_X1 \myidu/_1434_ ( .A(\myidu/_0484_ ), .B1(\myidu/_0535_ ), .B2(\myidu/_0543_ ), .ZN(\myidu/_0544_ ) );
NAND2_X1 \myidu/_1435_ ( .A1(\myidu/_0528_ ), .A2(\myidu/_0794_ ), .ZN(\myidu/_0545_ ) );
AOI21_X1 \myidu/_1436_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0544_ ), .B2(\myidu/_0545_ ), .ZN(\myidu/_0042_ ) );
NAND2_X1 \myidu/_1437_ ( .A1(\myidu/_0500_ ), .A2(\myidu/_0429_ ), .ZN(\myidu/_0546_ ) );
AND2_X1 \myidu/_1438_ ( .A1(\myidu/_0540_ ), .A2(\myidu/_0546_ ), .ZN(\myidu/_0547_ ) );
AND3_X1 \myidu/_1439_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0264_ ), .A3(\myidu/_0509_ ), .ZN(\myidu/_0548_ ) );
AOI21_X1 \myidu/_1440_ ( .A(\myidu/_0548_ ), .B1(\myidu/_0159_ ), .B2(\myidu/_0235_ ), .ZN(\myidu/_0549_ ) );
OAI21_X1 \myidu/_1441_ ( .A(\myidu/_0209_ ), .B1(\myidu/_0494_ ), .B2(\myidu/_0506_ ), .ZN(\myidu/_0550_ ) );
NAND4_X1 \myidu/_1442_ ( .A1(\myidu/_0547_ ), .A2(\myidu/_0377_ ), .A3(\myidu/_0549_ ), .A4(\myidu/_0550_ ), .ZN(\myidu/_0551_ ) );
NAND4_X1 \myidu/_1443_ ( .A1(\myidu/_0305_ ), .A2(\myidu/_0485_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0301_ ), .ZN(\myidu/_0552_ ) );
NAND4_X1 \myidu/_1444_ ( .A1(\myidu/_0293_ ), .A2(\myidu/_0485_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0301_ ), .ZN(\myidu/_0553_ ) );
AOI21_X1 \myidu/_1445_ ( .A(\myidu/_0179_ ), .B1(\myidu/_0552_ ), .B2(\myidu/_0553_ ), .ZN(\myidu/_0554_ ) );
NAND4_X1 \myidu/_1446_ ( .A1(\myidu/_0285_ ), .A2(\myidu/_0485_ ), .A3(\myidu/_0201_ ), .A4(\myidu/_0301_ ), .ZN(\myidu/_0555_ ) );
NOR2_X1 \myidu/_1447_ ( .A1(\myidu/_0555_ ), .A2(\myidu/_0179_ ), .ZN(\myidu/_0556_ ) );
NOR2_X1 \myidu/_1448_ ( .A1(\myidu/_0554_ ), .A2(\myidu/_0556_ ), .ZN(\myidu/_0557_ ) );
AOI21_X1 \myidu/_1449_ ( .A(\myidu/_0210_ ), .B1(\myidu/_0518_ ), .B2(\myidu/_0429_ ), .ZN(\myidu/_0558_ ) );
NAND2_X1 \myidu/_1450_ ( .A1(\myidu/_0557_ ), .A2(\myidu/_0558_ ), .ZN(\myidu/_0559_ ) );
OAI21_X1 \myidu/_1451_ ( .A(\myidu/_0484_ ), .B1(\myidu/_0551_ ), .B2(\myidu/_0559_ ), .ZN(\myidu/_0560_ ) );
NAND2_X1 \myidu/_1452_ ( .A1(\myidu/_0528_ ), .A2(\myidu/_0795_ ), .ZN(\myidu/_0561_ ) );
AOI21_X1 \myidu/_1453_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0560_ ), .B2(\myidu/_0561_ ), .ZN(\myidu/_0043_ ) );
AND2_X1 \myidu/_1454_ ( .A1(\myidu/_0273_ ), .A2(\myidu/_0287_ ), .ZN(\myidu/_0562_ ) );
AND4_X1 \myidu/_1455_ ( .A1(\myidu/_0486_ ), .A2(\myidu/_0562_ ), .A3(\myidu/_0302_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0563_ ) );
OAI21_X1 \myidu/_1456_ ( .A(\myidu/_0290_ ), .B1(\myidu/_0563_ ), .B2(\myidu/_0519_ ), .ZN(\myidu/_0564_ ) );
NAND4_X1 \myidu/_1457_ ( .A1(\myidu/_0343_ ), .A2(\myidu/_0176_ ), .A3(\myidu/_0175_ ), .A4(\myidu/_0344_ ), .ZN(\myidu/_0565_ ) );
NAND4_X1 \myidu/_1458_ ( .A1(\myidu/_0338_ ), .A2(\myidu/_0368_ ), .A3(\myidu/_0168_ ), .A4(\myidu/_0340_ ), .ZN(\myidu/_0566_ ) );
NOR2_X1 \myidu/_1459_ ( .A1(\myidu/_0565_ ), .A2(\myidu/_0566_ ), .ZN(\myidu/_0567_ ) );
NAND2_X1 \myidu/_1460_ ( .A1(\myidu/_0567_ ), .A2(\myidu/_0356_ ), .ZN(\myidu/_0568_ ) );
AND2_X1 \myidu/_1461_ ( .A1(\myidu/_0523_ ), .A2(\myidu/_0209_ ), .ZN(\myidu/_0569_ ) );
NOR2_X1 \myidu/_1462_ ( .A1(\myidu/_0569_ ), .A2(\myidu/_0376_ ), .ZN(\myidu/_0570_ ) );
NAND4_X1 \myidu/_1463_ ( .A1(\myidu/_0564_ ), .A2(\myidu/_0495_ ), .A3(\myidu/_0568_ ), .A4(\myidu/_0570_ ), .ZN(\myidu/_0571_ ) );
MUX2_X1 \myidu/_1464_ ( .A(\myidu/_0796_ ), .B(\myidu/_0571_ ), .S(\myidu/_0320_ ), .Z(\myidu/_0572_ ) );
AND2_X1 \myidu/_1465_ ( .A1(\myidu/_0572_ ), .A2(\myidu/_0325_ ), .ZN(\myidu/_0044_ ) );
BUF_X4 \myidu/_1466_ ( .A(\myidu/_0323_ ), .Z(\myidu/_0573_ ) );
OAI21_X1 \myidu/_1467_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0320_ ), .B2(\myidu/_0797_ ), .ZN(\myidu/_0574_ ) );
NAND2_X1 \myidu/_1468_ ( .A1(\myidu/_0295_ ), .A2(\myidu/_0570_ ), .ZN(\myidu/_0575_ ) );
NAND2_X1 \myidu/_1469_ ( .A1(\myidu/_0213_ ), .A2(\myidu/_0228_ ), .ZN(\myidu/_0576_ ) );
AND2_X1 \myidu/_1470_ ( .A1(\myidu/_0576_ ), .A2(\myidu/_0225_ ), .ZN(\myidu/_0577_ ) );
INV_X1 \myidu/_1471_ ( .A(\myidu/_0577_ ), .ZN(\myidu/_0578_ ) );
NOR3_X1 \myidu/_1472_ ( .A1(\myidu/_0575_ ), .A2(\myidu/_0362_ ), .A3(\myidu/_0578_ ), .ZN(\myidu/_0579_ ) );
AOI21_X1 \myidu/_1473_ ( .A(\myidu/_0574_ ), .B1(\myidu/_0579_ ), .B2(\myidu/_0484_ ), .ZN(\myidu/_0045_ ) );
NAND4_X1 \myidu/_1474_ ( .A1(\myidu/_0285_ ), .A2(\myidu/_0485_ ), .A3(\myidu/_0301_ ), .A4(\myidu/_0212_ ), .ZN(\myidu/_0580_ ) );
NOR2_X1 \myidu/_1475_ ( .A1(\myidu/_0580_ ), .A2(\myidu/_0179_ ), .ZN(\myidu/_0581_ ) );
NAND4_X1 \myidu/_1476_ ( .A1(\myidu/_0517_ ), .A2(\myidu/_0485_ ), .A3(\myidu/_0201_ ), .A4(\myidu/_0300_ ), .ZN(\myidu/_0582_ ) );
NAND4_X1 \myidu/_1477_ ( .A1(\myidu/_0562_ ), .A2(\myidu/_0211_ ), .A3(\myidu/_0300_ ), .A4(\myidu/_0212_ ), .ZN(\myidu/_0583_ ) );
AOI21_X1 \myidu/_1478_ ( .A(\myidu/_0179_ ), .B1(\myidu/_0582_ ), .B2(\myidu/_0583_ ), .ZN(\myidu/_0584_ ) );
AOI211_X4 \myidu/_1479_ ( .A(\myidu/_0581_ ), .B(\myidu/_0584_ ), .C1(\myidu/_0360_ ), .C2(\myidu/_0523_ ), .ZN(\myidu/_0585_ ) );
NAND4_X1 \myidu/_1480_ ( .A1(\myidu/_0299_ ), .A2(\myidu/_0297_ ), .A3(\myidu/_0308_ ), .A4(\myidu/_0301_ ), .ZN(\myidu/_0586_ ) );
NAND4_X1 \myidu/_1481_ ( .A1(\myidu/_0299_ ), .A2(\myidu/_0297_ ), .A3(\myidu/_0301_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0587_ ) );
AOI21_X1 \myidu/_1482_ ( .A(\myidu/_0179_ ), .B1(\myidu/_0586_ ), .B2(\myidu/_0587_ ), .ZN(\myidu/_0588_ ) );
NAND4_X1 \myidu/_1483_ ( .A1(\myidu/_0305_ ), .A2(\myidu/_0485_ ), .A3(\myidu/_0301_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0589_ ) );
AOI21_X1 \myidu/_1484_ ( .A(\myidu/_0179_ ), .B1(\myidu/_0589_ ), .B2(\myidu/_0555_ ), .ZN(\myidu/_0590_ ) );
NAND4_X1 \myidu/_1485_ ( .A1(\myidu/_0293_ ), .A2(\myidu/_0297_ ), .A3(\myidu/_0301_ ), .A4(\myidu/_0303_ ), .ZN(\myidu/_0591_ ) );
NOR2_X1 \myidu/_1486_ ( .A1(\myidu/_0591_ ), .A2(\myidu/_0179_ ), .ZN(\myidu/_0592_ ) );
NOR4_X1 \myidu/_1487_ ( .A1(\myidu/_0588_ ), .A2(\myidu/_0554_ ), .A3(\myidu/_0590_ ), .A4(\myidu/_0592_ ), .ZN(\myidu/_0593_ ) );
OAI21_X1 \myidu/_1488_ ( .A(\myidu/_0221_ ), .B1(\myidu/_0207_ ), .B2(\myidu/_0523_ ), .ZN(\myidu/_0594_ ) );
AOI22_X1 \myidu/_1489_ ( .A1(\myidu/_0207_ ), .A2(\myidu/_0209_ ), .B1(\myidu/_0489_ ), .B2(\myidu/_0523_ ), .ZN(\myidu/_0595_ ) );
NAND4_X1 \myidu/_1490_ ( .A1(\myidu/_0585_ ), .A2(\myidu/_0593_ ), .A3(\myidu/_0594_ ), .A4(\myidu/_0595_ ), .ZN(\myidu/_0596_ ) );
NAND2_X1 \myidu/_1491_ ( .A1(\myidu/_0506_ ), .A2(\myidu/_0209_ ), .ZN(\myidu/_0597_ ) );
AND2_X1 \myidu/_1492_ ( .A1(\myidu/_0597_ ), .A2(\myidu/_0536_ ), .ZN(\myidu/_0598_ ) );
NAND2_X1 \myidu/_1493_ ( .A1(\myidu/_0506_ ), .A2(\myidu/_0360_ ), .ZN(\myidu/_0599_ ) );
NAND4_X1 \myidu/_1494_ ( .A1(\myidu/_0598_ ), .A2(\myidu/_0599_ ), .A3(\myidu/_0507_ ), .A4(\myidu/_0537_ ), .ZN(\myidu/_0600_ ) );
NAND2_X1 \myidu/_1495_ ( .A1(\myidu/_0370_ ), .A2(\myidu/_0356_ ), .ZN(\myidu/_0601_ ) );
NAND3_X1 \myidu/_1496_ ( .A1(\myidu/_0601_ ), .A2(\myidu/_0493_ ), .A3(\myidu/_0392_ ), .ZN(\myidu/_0602_ ) );
OR4_X1 \myidu/_1497_ ( .A1(\myidu/_0575_ ), .A2(\myidu/_0596_ ), .A3(\myidu/_0600_ ), .A4(\myidu/_0602_ ), .ZN(\myidu/_0603_ ) );
MUX2_X1 \myidu/_1498_ ( .A(\myidu/_0798_ ), .B(\myidu/_0603_ ), .S(\myidu/_0320_ ), .Z(\myidu/_0604_ ) );
AND2_X1 \myidu/_1499_ ( .A1(\myidu/_0604_ ), .A2(\myidu/_0325_ ), .ZN(\myidu/_0046_ ) );
AND2_X1 \myidu/_1500_ ( .A1(\myidu/_0370_ ), .A2(\myidu/_0366_ ), .ZN(\myidu/_0605_ ) );
NOR2_X1 \myidu/_1501_ ( .A1(\myidu/_0605_ ), .A2(\myidu/_0332_ ), .ZN(\myidu/_0606_ ) );
INV_X1 \myidu/_1502_ ( .A(\myidu/_0606_ ), .ZN(\myidu/_0607_ ) );
AOI21_X1 \myidu/_1503_ ( .A(\myidu/_0498_ ), .B1(\myidu/_0494_ ), .B2(\myidu/_0360_ ), .ZN(\myidu/_0608_ ) );
AND3_X1 \myidu/_1504_ ( .A1(\myidu/_0216_ ), .A2(\myidu/_0486_ ), .A3(\myidu/_0360_ ), .ZN(\myidu/_0609_ ) );
AOI21_X1 \myidu/_1505_ ( .A(\myidu/_0609_ ), .B1(\myidu/_0489_ ), .B2(\myidu/_0506_ ), .ZN(\myidu/_0610_ ) );
AOI22_X1 \myidu/_1506_ ( .A1(\myidu/_0209_ ), .A2(\myidu/_0494_ ), .B1(\myidu/_0506_ ), .B2(\myidu/_0360_ ), .ZN(\myidu/_0611_ ) );
NAND4_X1 \myidu/_1507_ ( .A1(\myidu/_0598_ ), .A2(\myidu/_0608_ ), .A3(\myidu/_0610_ ), .A4(\myidu/_0611_ ), .ZN(\myidu/_0612_ ) );
OAI21_X1 \myidu/_1508_ ( .A(\myidu/_0484_ ), .B1(\myidu/_0607_ ), .B2(\myidu/_0612_ ), .ZN(\myidu/_0613_ ) );
NAND2_X1 \myidu/_1509_ ( .A1(\myidu/_0528_ ), .A2(\myidu/_0799_ ), .ZN(\myidu/_0614_ ) );
AOI21_X1 \myidu/_1510_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0613_ ), .B2(\myidu/_0614_ ), .ZN(\myidu/_0047_ ) );
AOI22_X1 \myidu/_1511_ ( .A1(\myidu/_0183_ ), .A2(\myidu/_0266_ ), .B1(\myidu/_0373_ ), .B2(\myidu/_0366_ ), .ZN(\myidu/_0615_ ) );
NOR2_X1 \myidu/_1512_ ( .A1(\myidu/_0199_ ), .A2(\myidu/_0391_ ), .ZN(\myidu/_0616_ ) );
AND4_X1 \myidu/_1513_ ( .A1(\myidu/_0319_ ), .A2(\myidu/_0615_ ), .A3(\myidu/_0483_ ), .A4(\myidu/_0616_ ), .ZN(\myidu/_0617_ ) );
AOI221_X4 \myidu/_1514_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0246_ ), .B2(\myidu/_0527_ ), .C1(\myidu/_0617_ ), .C2(\myidu/_0606_ ), .ZN(\myidu/_0048_ ) );
BUF_X4 \myidu/_1515_ ( .A(\myidu/_0400_ ), .Z(\myidu/_0618_ ) );
OAI21_X1 \myidu/_1516_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0779_ ), .ZN(\myidu/_0619_ ) );
BUF_X4 \myidu/_1517_ ( .A(\myidu/_0400_ ), .Z(\myidu/_0620_ ) );
AND2_X2 \myidu/_1518_ ( .A1(\myidu/_0363_ ), .A2(\myidu/_0374_ ), .ZN(\myidu/_0621_ ) );
NAND3_X1 \myidu/_1519_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0161_ ), .A3(\myidu/_0434_ ), .ZN(\myidu/_0622_ ) );
AOI21_X1 \myidu/_1520_ ( .A(\myidu/_0619_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0622_ ), .ZN(\myidu/_0081_ ) );
OAI21_X1 \myidu/_1521_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0780_ ), .ZN(\myidu/_0623_ ) );
NAND3_X1 \myidu/_1522_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0162_ ), .A3(\myidu/_0434_ ), .ZN(\myidu/_0624_ ) );
AOI21_X1 \myidu/_1523_ ( .A(\myidu/_0623_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0624_ ), .ZN(\myidu/_0082_ ) );
OAI21_X1 \myidu/_1524_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0781_ ), .ZN(\myidu/_0625_ ) );
NAND3_X1 \myidu/_1525_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0163_ ), .A3(\myidu/_0434_ ), .ZN(\myidu/_0626_ ) );
AOI21_X1 \myidu/_1526_ ( .A(\myidu/_0625_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0626_ ), .ZN(\myidu/_0083_ ) );
INV_X1 \myidu/_1527_ ( .A(\myidu/_0400_ ), .ZN(\myidu/_0627_ ) );
AND2_X1 \myidu/_1528_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0434_ ), .ZN(\myidu/_0628_ ) );
AOI21_X1 \myidu/_1529_ ( .A(\myidu/_0627_ ), .B1(\myidu/_0164_ ), .B2(\myidu/_0628_ ), .ZN(\myidu/_0629_ ) );
OAI21_X1 \myidu/_1530_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0782_ ), .ZN(\myidu/_0630_ ) );
NOR2_X1 \myidu/_1531_ ( .A1(\myidu/_0629_ ), .A2(\myidu/_0630_ ), .ZN(\myidu/_0084_ ) );
OAI21_X1 \myidu/_1532_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0783_ ), .ZN(\myidu/_0631_ ) );
NAND3_X1 \myidu/_1533_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0165_ ), .A3(\myidu/_0434_ ), .ZN(\myidu/_0632_ ) );
AOI21_X1 \myidu/_1534_ ( .A(\myidu/_0631_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0632_ ), .ZN(\myidu/_0085_ ) );
NAND2_X1 \myidu/_1535_ ( .A1(\myidu/_0207_ ), .A2(\myidu/_0221_ ), .ZN(\myidu/_0633_ ) );
NAND2_X1 \myidu/_1536_ ( .A1(\myidu/_0633_ ), .A2(\myidu/_0576_ ), .ZN(\myidu/_0634_ ) );
AND2_X1 \myidu/_1537_ ( .A1(\myidu/_0373_ ), .A2(\myidu/_0366_ ), .ZN(\myidu/_0635_ ) );
NOR4_X1 \myidu/_1538_ ( .A1(\myidu/_0607_ ), .A2(\myidu/_0634_ ), .A3(\myidu/_0635_ ), .A4(\myidu/_0575_ ), .ZN(\myidu/_0636_ ) );
NAND3_X1 \myidu/_1539_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0360_ ), .A3(\myidu/_0215_ ), .ZN(\myidu/_0637_ ) );
AND4_X1 \myidu/_1540_ ( .A1(\myidu/_0220_ ), .A2(\myidu/_0364_ ), .A3(\myidu/_0222_ ), .A4(\myidu/_0215_ ), .ZN(\myidu/_0638_ ) );
NOR3_X1 \myidu/_1541_ ( .A1(\myidu/_0210_ ), .A2(\myidu/_0638_ ), .A3(\myidu/_0218_ ), .ZN(\myidu/_0639_ ) );
AND4_X1 \myidu/_1542_ ( .A1(\myidu/_0637_ ), .A2(\myidu/_0363_ ), .A3(\myidu/_0616_ ), .A4(\myidu/_0639_ ), .ZN(\myidu/_0640_ ) );
AND2_X1 \myidu/_1543_ ( .A1(\myidu/_0636_ ), .A2(\myidu/_0640_ ), .ZN(\myidu/_0641_ ) );
AOI211_X4 \myidu/_1544_ ( .A(\myidu/_0527_ ), .B(\myidu/_0398_ ), .C1(\myidu/_0641_ ), .C2(\myidu/_0167_ ), .ZN(\myidu/_0642_ ) );
OAI21_X1 \myidu/_1545_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0784_ ), .ZN(\myidu/_0643_ ) );
NOR2_X1 \myidu/_1546_ ( .A1(\myidu/_0642_ ), .A2(\myidu/_0643_ ), .ZN(\myidu/_0086_ ) );
AOI211_X4 \myidu/_1547_ ( .A(\myidu/_0527_ ), .B(\myidu/_0398_ ), .C1(\myidu/_0641_ ), .C2(\myidu/_0168_ ), .ZN(\myidu/_0644_ ) );
OAI21_X1 \myidu/_1548_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0785_ ), .ZN(\myidu/_0645_ ) );
NOR2_X1 \myidu/_1549_ ( .A1(\myidu/_0644_ ), .A2(\myidu/_0645_ ), .ZN(\myidu/_0087_ ) );
AOI211_X4 \myidu/_1550_ ( .A(\myidu/_0527_ ), .B(\myidu/_0398_ ), .C1(\myidu/_0641_ ), .C2(\myidu/_0169_ ), .ZN(\myidu/_0646_ ) );
OAI21_X1 \myidu/_1551_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0786_ ), .ZN(\myidu/_0647_ ) );
NOR2_X1 \myidu/_1552_ ( .A1(\myidu/_0646_ ), .A2(\myidu/_0647_ ), .ZN(\myidu/_0088_ ) );
AOI211_X4 \myidu/_1553_ ( .A(\myidu/_0527_ ), .B(\myidu/_0398_ ), .C1(\myidu/_0641_ ), .C2(\myidu/_0170_ ), .ZN(\myidu/_0648_ ) );
OAI21_X1 \myidu/_1554_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0787_ ), .ZN(\myidu/_0649_ ) );
NOR2_X1 \myidu/_1555_ ( .A1(\myidu/_0648_ ), .A2(\myidu/_0649_ ), .ZN(\myidu/_0089_ ) );
AOI211_X4 \myidu/_1556_ ( .A(\myidu/_0527_ ), .B(\myidu/_0398_ ), .C1(\myidu/_0641_ ), .C2(\myidu/_0171_ ), .ZN(\myidu/_0650_ ) );
OAI21_X1 \myidu/_1557_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0788_ ), .ZN(\myidu/_0651_ ) );
NOR2_X1 \myidu/_1558_ ( .A1(\myidu/_0650_ ), .A2(\myidu/_0651_ ), .ZN(\myidu/_0090_ ) );
AND2_X1 \myidu/_1559_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0268_ ), .ZN(\myidu/_0652_ ) );
AOI21_X1 \myidu/_1560_ ( .A(\myidu/_0627_ ), .B1(\myidu/_0184_ ), .B2(\myidu/_0652_ ), .ZN(\myidu/_0653_ ) );
OAI21_X1 \myidu/_1561_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0772_ ), .ZN(\myidu/_0654_ ) );
NOR2_X1 \myidu/_1562_ ( .A1(\myidu/_0653_ ), .A2(\myidu/_0654_ ), .ZN(\myidu/_0091_ ) );
OAI21_X1 \myidu/_1563_ ( .A(\myidu/_0323_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0773_ ), .ZN(\myidu/_0655_ ) );
NAND3_X1 \myidu/_1564_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0185_ ), .A3(\myidu/_0268_ ), .ZN(\myidu/_0656_ ) );
AOI21_X1 \myidu/_1565_ ( .A(\myidu/_0655_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0656_ ), .ZN(\myidu/_0092_ ) );
AOI21_X1 \myidu/_1566_ ( .A(\myidu/_0627_ ), .B1(\myidu/_0186_ ), .B2(\myidu/_0652_ ), .ZN(\myidu/_0657_ ) );
OAI21_X1 \myidu/_1567_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0774_ ), .ZN(\myidu/_0658_ ) );
NOR2_X1 \myidu/_1568_ ( .A1(\myidu/_0657_ ), .A2(\myidu/_0658_ ), .ZN(\myidu/_0093_ ) );
AOI21_X1 \myidu/_1569_ ( .A(\myidu/_0627_ ), .B1(\myidu/_0156_ ), .B2(\myidu/_0652_ ), .ZN(\myidu/_0659_ ) );
OAI21_X1 \myidu/_1570_ ( .A(\myidu/_0573_ ), .B1(\myidu/_0618_ ), .B2(\myidu/_0775_ ), .ZN(\myidu/_0660_ ) );
NOR2_X1 \myidu/_1571_ ( .A1(\myidu/_0659_ ), .A2(\myidu/_0660_ ), .ZN(\myidu/_0094_ ) );
OAI21_X1 \myidu/_1572_ ( .A(\myidu/_0323_ ), .B1(\myidu/_0400_ ), .B2(\myidu/_0776_ ), .ZN(\myidu/_0661_ ) );
NAND3_X1 \myidu/_1573_ ( .A1(\myidu/_0621_ ), .A2(\myidu/_0157_ ), .A3(\myidu/_0268_ ), .ZN(\myidu/_0662_ ) );
AOI21_X1 \myidu/_1574_ ( .A(\myidu/_0661_ ), .B1(\myidu/_0620_ ), .B2(\myidu/_0662_ ), .ZN(\myidu/_0095_ ) );
INV_X1 \myidu/_1575_ ( .A(\myidu/_0635_ ), .ZN(\myidu/_0663_ ) );
AND2_X2 \myidu/_1576_ ( .A1(\myidu/_0606_ ), .A2(\myidu/_0663_ ), .ZN(\myidu/_0664_ ) );
NOR2_X1 \myidu/_1577_ ( .A1(\myidu/_0664_ ), .A2(\myidu/_0527_ ), .ZN(\myidu/_0665_ ) );
OAI21_X1 \myidu/_1578_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0110_ ), .ZN(\myidu/_0666_ ) );
NAND3_X1 \myidu/_1579_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0368_ ), .A3(\myidu/_0320_ ), .ZN(\myidu/_0667_ ) );
INV_X1 \myidu/_1580_ ( .A(\myidu/_0667_ ), .ZN(\myidu/_0668_ ) );
NOR2_X1 \myidu/_1581_ ( .A1(\myidu/_0666_ ), .A2(\myidu/_0668_ ), .ZN(\myidu/_0096_ ) );
OAI21_X1 \myidu/_1582_ ( .A(\myidu/_0113_ ), .B1(\myidu/_0664_ ), .B2(\myidu/_0528_ ), .ZN(\myidu/_0669_ ) );
NAND3_X1 \myidu/_1583_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0168_ ), .A3(\myidu/_0484_ ), .ZN(\myidu/_0670_ ) );
AOI21_X1 \myidu/_1584_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0669_ ), .B2(\myidu/_0670_ ), .ZN(\myidu/_0097_ ) );
OAI21_X1 \myidu/_1585_ ( .A(\myidu/_0323_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0114_ ), .ZN(\myidu/_0671_ ) );
AND2_X1 \myidu/_1586_ ( .A1(\myidu/_0370_ ), .A2(\myidu/_0356_ ), .ZN(\myidu/_0672_ ) );
AOI21_X1 \myidu/_1587_ ( .A(\myidu/_0672_ ), .B1(\myidu/_0169_ ), .B2(\myidu/_0333_ ), .ZN(\myidu/_0673_ ) );
AOI21_X1 \myidu/_1588_ ( .A(\myidu/_0671_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0673_ ), .ZN(\myidu/_0098_ ) );
OAI21_X1 \myidu/_1589_ ( .A(\myidu/_0115_ ), .B1(\myidu/_0664_ ), .B2(\myidu/_0528_ ), .ZN(\myidu/_0674_ ) );
NAND3_X1 \myidu/_1590_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0170_ ), .A3(\myidu/_0484_ ), .ZN(\myidu/_0675_ ) );
AOI21_X1 \myidu/_1591_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0674_ ), .B2(\myidu/_0675_ ), .ZN(\myidu/_0099_ ) );
OAI21_X1 \myidu/_1592_ ( .A(\myidu/_0116_ ), .B1(\myidu/_0664_ ), .B2(\myidu/_0528_ ), .ZN(\myidu/_0676_ ) );
NAND3_X1 \myidu/_1593_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0171_ ), .A3(\myidu/_0484_ ), .ZN(\myidu/_0677_ ) );
AOI21_X1 \myidu/_1594_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0676_ ), .B2(\myidu/_0677_ ), .ZN(\myidu/_0100_ ) );
OAI21_X1 \myidu/_1595_ ( .A(\myidu/_0117_ ), .B1(\myidu/_0664_ ), .B2(\myidu/_0528_ ), .ZN(\myidu/_0678_ ) );
NAND3_X1 \myidu/_1596_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0172_ ), .A3(\myidu/_0484_ ), .ZN(\myidu/_0679_ ) );
AOI21_X1 \myidu/_1597_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0678_ ), .B2(\myidu/_0679_ ), .ZN(\myidu/_0101_ ) );
OAI21_X1 \myidu/_1598_ ( .A(\myidu/_0323_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0118_ ), .ZN(\myidu/_0680_ ) );
MUX2_X1 \myidu/_1599_ ( .A(\myidu/_0283_ ), .B(\myidu/_0605_ ), .S(\myidu/_0236_ ), .Z(\myidu/_0681_ ) );
AOI21_X1 \myidu/_1600_ ( .A(\myidu/_0680_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0681_ ), .ZN(\myidu/_0102_ ) );
OAI221_X1 \myidu/_1601_ ( .A(\myidu/_0320_ ), .B1(\myidu/_0272_ ), .B2(\myidu/_0236_ ), .C1(\myidu/_0607_ ), .C2(\myidu/_0635_ ), .ZN(\myidu/_0682_ ) );
OAI21_X1 \myidu/_1602_ ( .A(\myidu/_0682_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0119_ ), .ZN(\myidu/_0683_ ) );
NOR2_X1 \myidu/_1603_ ( .A1(\myidu/_0683_ ), .A2(\myidu/_0789_ ), .ZN(\myidu/_0103_ ) );
OAI21_X1 \myidu/_1604_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0120_ ), .ZN(\myidu/_0684_ ) );
OR3_X1 \myidu/_1605_ ( .A1(\myidu/_0236_ ), .A2(\myidu/_0175_ ), .A3(\myidu/_0527_ ), .ZN(\myidu/_0685_ ) );
INV_X1 \myidu/_1606_ ( .A(\myidu/_0685_ ), .ZN(\myidu/_0686_ ) );
NOR2_X1 \myidu/_1607_ ( .A1(\myidu/_0684_ ), .A2(\myidu/_0686_ ), .ZN(\myidu/_0104_ ) );
OAI21_X1 \myidu/_1608_ ( .A(\myidu/_0325_ ), .B1(\myidu/_0665_ ), .B2(\myidu/_0121_ ), .ZN(\myidu/_0687_ ) );
OR3_X1 \myidu/_1609_ ( .A1(\myidu/_0236_ ), .A2(\myidu/_0176_ ), .A3(\myidu/_0527_ ), .ZN(\myidu/_0688_ ) );
INV_X1 \myidu/_1610_ ( .A(\myidu/_0688_ ), .ZN(\myidu/_0689_ ) );
NOR2_X1 \myidu/_1611_ ( .A1(\myidu/_0687_ ), .A2(\myidu/_0689_ ), .ZN(\myidu/_0105_ ) );
OAI21_X1 \myidu/_1612_ ( .A(\myidu/_0111_ ), .B1(\myidu/_0664_ ), .B2(\myidu/_0528_ ), .ZN(\myidu/_0690_ ) );
NAND3_X1 \myidu/_1613_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0178_ ), .A3(\myidu/_0320_ ), .ZN(\myidu/_0691_ ) );
AOI21_X1 \myidu/_1614_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0690_ ), .B2(\myidu/_0691_ ), .ZN(\myidu/_0106_ ) );
OAI21_X1 \myidu/_1615_ ( .A(\myidu/_0112_ ), .B1(\myidu/_0664_ ), .B2(\myidu/_0528_ ), .ZN(\myidu/_0692_ ) );
NAND3_X1 \myidu/_1616_ ( .A1(\myidu/_0333_ ), .A2(\myidu/_0179_ ), .A3(\myidu/_0320_ ), .ZN(\myidu/_0693_ ) );
AOI21_X1 \myidu/_1617_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0692_ ), .B2(\myidu/_0693_ ), .ZN(\myidu/_0107_ ) );
AND2_X1 \myidu/_1618_ ( .A1(\myidu/_0238_ ), .A2(\myidu/_0249_ ), .ZN(\myidu/_0694_ ) );
AND3_X1 \myidu/_1619_ ( .A1(\myidu/_0237_ ), .A2(\myidu/_0258_ ), .A3(\myidu/_0628_ ), .ZN(\myidu/_0695_ ) );
OAI21_X1 \myidu/_1620_ ( .A(\myidu/_0778_ ), .B1(\myidu/_0694_ ), .B2(\myidu/_0695_ ), .ZN(\myidu/_0696_ ) );
AND2_X1 \myidu/_1621_ ( .A1(\myidu/_0237_ ), .A2(\myidu/_0628_ ), .ZN(\myidu/_0697_ ) );
INV_X1 \myidu/_1622_ ( .A(\myidu/_0007_ ), .ZN(\myidu/_0698_ ) );
NOR2_X1 \myidu/_1623_ ( .A1(\myidu/_0296_ ), .A2(\myidu/_0386_ ), .ZN(\myidu/_0699_ ) );
AND3_X2 \myidu/_1624_ ( .A1(\myidu/_0697_ ), .A2(\myidu/_0698_ ), .A3(\myidu/_0699_ ), .ZN(\myidu/_0700_ ) );
NOR2_X1 \myidu/_1625_ ( .A1(\myidu/_0329_ ), .A2(\myidu/_0187_ ), .ZN(\myidu/_0701_ ) );
NOR3_X1 \myidu/_1626_ ( .A1(\myidu/_0189_ ), .A2(\myidu/_0481_ ), .A3(\myidu/_0701_ ), .ZN(\myidu/_0702_ ) );
INV_X1 \myidu/_1627_ ( .A(\myidu/_0702_ ), .ZN(\myidu/_0703_ ) );
OR3_X1 \myidu/_1628_ ( .A1(\myidu/_0696_ ), .A2(\myidu/_0700_ ), .A3(\myidu/_0703_ ), .ZN(\myidu/_0704_ ) );
OAI21_X1 \myidu/_1629_ ( .A(\myidu/_0791_ ), .B1(\myidu/_0700_ ), .B2(\myidu/_0703_ ), .ZN(\myidu/_0705_ ) );
AOI21_X1 \myidu/_1630_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0704_ ), .B2(\myidu/_0705_ ), .ZN(\myidu/_0108_ ) );
OAI21_X1 \myidu/_1631_ ( .A(\myidu/_0122_ ), .B1(\myidu/_0189_ ), .B2(\myidu/_0698_ ), .ZN(\myidu/_0706_ ) );
OAI211_X2 \myidu/_1632_ ( .A(\myidu/_0792_ ), .B(\myidu/_0007_ ), .C1(\myidu/_0188_ ), .C2(\myidu/_0777_ ), .ZN(\myidu/_0707_ ) );
AOI21_X1 \myidu/_1633_ ( .A(\myidu/_0789_ ), .B1(\myidu/_0706_ ), .B2(\myidu/_0707_ ), .ZN(\myidu/_0109_ ) );
DFF_X1 \myidu/_1634_ ( .D(\myidu/_0000_ ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu/_0003_ ) );
DFF_X1 \myidu/_1635_ ( .D(\myidu/_0001_ ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu/_0906_ ) );
DFF_X1 \myidu/_1636_ ( .D(\myidu/_0002_ ), .CK(clock ), .Q(\myidu/state [2] ), .QN(\myidu/_0905_ ) );
DFF_X1 \myidu/_1637_ ( .D(\myidu/_0907_ ), .CK(clock ), .Q(\ID_EX_imm [0] ), .QN(\myidu/_0904_ ) );
DFF_X1 \myidu/_1638_ ( .D(\myidu/_0908_ ), .CK(clock ), .Q(\ID_EX_imm [1] ), .QN(\myidu/_0903_ ) );
DFF_X1 \myidu/_1639_ ( .D(\myidu/_0909_ ), .CK(clock ), .Q(\ID_EX_imm [2] ), .QN(\myidu/_0902_ ) );
DFF_X1 \myidu/_1640_ ( .D(\myidu/_0910_ ), .CK(clock ), .Q(\ID_EX_imm [3] ), .QN(\myidu/_0901_ ) );
DFF_X1 \myidu/_1641_ ( .D(\myidu/_0911_ ), .CK(clock ), .Q(\ID_EX_imm [4] ), .QN(\myidu/_0900_ ) );
DFF_X1 \myidu/_1642_ ( .D(\myidu/_0912_ ), .CK(clock ), .Q(\ID_EX_imm [5] ), .QN(\myidu/_0899_ ) );
DFF_X1 \myidu/_1643_ ( .D(\myidu/_0913_ ), .CK(clock ), .Q(\ID_EX_imm [6] ), .QN(\myidu/_0898_ ) );
DFF_X1 \myidu/_1644_ ( .D(\myidu/_0914_ ), .CK(clock ), .Q(\ID_EX_imm [7] ), .QN(\myidu/_0897_ ) );
DFF_X1 \myidu/_1645_ ( .D(\myidu/_0915_ ), .CK(clock ), .Q(\ID_EX_imm [8] ), .QN(\myidu/_0896_ ) );
DFF_X1 \myidu/_1646_ ( .D(\myidu/_0916_ ), .CK(clock ), .Q(\ID_EX_imm [9] ), .QN(\myidu/_0895_ ) );
DFF_X1 \myidu/_1647_ ( .D(\myidu/_0917_ ), .CK(clock ), .Q(\ID_EX_imm [10] ), .QN(\myidu/_0894_ ) );
DFF_X1 \myidu/_1648_ ( .D(\myidu/_0918_ ), .CK(clock ), .Q(\ID_EX_imm [11] ), .QN(\myidu/_0893_ ) );
DFF_X1 \myidu/_1649_ ( .D(\myidu/_0919_ ), .CK(clock ), .Q(\ID_EX_imm [12] ), .QN(\myidu/_0892_ ) );
DFF_X1 \myidu/_1650_ ( .D(\myidu/_0920_ ), .CK(clock ), .Q(\ID_EX_imm [13] ), .QN(\myidu/_0891_ ) );
DFF_X1 \myidu/_1651_ ( .D(\myidu/_0921_ ), .CK(clock ), .Q(\ID_EX_imm [14] ), .QN(\myidu/_0890_ ) );
DFF_X1 \myidu/_1652_ ( .D(\myidu/_0922_ ), .CK(clock ), .Q(\ID_EX_imm [15] ), .QN(\myidu/_0889_ ) );
DFF_X1 \myidu/_1653_ ( .D(\myidu/_0923_ ), .CK(clock ), .Q(\ID_EX_imm [16] ), .QN(\myidu/_0888_ ) );
DFF_X1 \myidu/_1654_ ( .D(\myidu/_0924_ ), .CK(clock ), .Q(\ID_EX_imm [17] ), .QN(\myidu/_0887_ ) );
DFF_X1 \myidu/_1655_ ( .D(\myidu/_0925_ ), .CK(clock ), .Q(\ID_EX_imm [18] ), .QN(\myidu/_0886_ ) );
DFF_X1 \myidu/_1656_ ( .D(\myidu/_0926_ ), .CK(clock ), .Q(\ID_EX_imm [19] ), .QN(\myidu/_0885_ ) );
DFF_X1 \myidu/_1657_ ( .D(\myidu/_0927_ ), .CK(clock ), .Q(\ID_EX_imm [20] ), .QN(\myidu/_0884_ ) );
DFF_X1 \myidu/_1658_ ( .D(\myidu/_0928_ ), .CK(clock ), .Q(\ID_EX_imm [21] ), .QN(\myidu/_0883_ ) );
DFF_X1 \myidu/_1659_ ( .D(\myidu/_0929_ ), .CK(clock ), .Q(\ID_EX_imm [22] ), .QN(\myidu/_0882_ ) );
DFF_X1 \myidu/_1660_ ( .D(\myidu/_0930_ ), .CK(clock ), .Q(\ID_EX_imm [23] ), .QN(\myidu/_0881_ ) );
DFF_X1 \myidu/_1661_ ( .D(\myidu/_0931_ ), .CK(clock ), .Q(\ID_EX_imm [24] ), .QN(\myidu/_0880_ ) );
DFF_X1 \myidu/_1662_ ( .D(\myidu/_0932_ ), .CK(clock ), .Q(\ID_EX_imm [25] ), .QN(\myidu/_0879_ ) );
DFF_X1 \myidu/_1663_ ( .D(\myidu/_0933_ ), .CK(clock ), .Q(\ID_EX_imm [26] ), .QN(\myidu/_0878_ ) );
DFF_X1 \myidu/_1664_ ( .D(\myidu/_0934_ ), .CK(clock ), .Q(\ID_EX_imm [27] ), .QN(\myidu/_0877_ ) );
DFF_X1 \myidu/_1665_ ( .D(\myidu/_0935_ ), .CK(clock ), .Q(\ID_EX_imm [28] ), .QN(\myidu/_0876_ ) );
DFF_X1 \myidu/_1666_ ( .D(\myidu/_0936_ ), .CK(clock ), .Q(\ID_EX_imm [29] ), .QN(\myidu/_0875_ ) );
DFF_X1 \myidu/_1667_ ( .D(\myidu/_0937_ ), .CK(clock ), .Q(\ID_EX_imm [30] ), .QN(\myidu/_0874_ ) );
DFF_X1 \myidu/_1668_ ( .D(\myidu/_0938_ ), .CK(clock ), .Q(\ID_EX_imm [31] ), .QN(\myidu/_0873_ ) );
DFF_X1 \myidu/_1669_ ( .D(\myidu/_0939_ ), .CK(clock ), .Q(stall_quest_fencei ), .QN(\myidu/_0872_ ) );
DFF_X1 \myidu/_1670_ ( .D(\myidu/_0940_ ), .CK(clock ), .Q(\ID_EX_typ [0] ), .QN(\myidu/_0871_ ) );
DFF_X1 \myidu/_1671_ ( .D(\myidu/_0941_ ), .CK(clock ), .Q(\ID_EX_typ [1] ), .QN(\myidu/_0870_ ) );
DFF_X1 \myidu/_1672_ ( .D(\myidu/_0942_ ), .CK(clock ), .Q(\ID_EX_typ [2] ), .QN(\myidu/_0869_ ) );
DFF_X1 \myidu/_1673_ ( .D(\myidu/_0943_ ), .CK(clock ), .Q(\ID_EX_typ [3] ), .QN(\myidu/_0868_ ) );
DFF_X1 \myidu/_1674_ ( .D(\myidu/_0944_ ), .CK(clock ), .Q(\ID_EX_typ [4] ), .QN(\myidu/_0867_ ) );
DFF_X1 \myidu/_1675_ ( .D(\myidu/_0945_ ), .CK(clock ), .Q(\ID_EX_typ [5] ), .QN(\myidu/_0866_ ) );
DFF_X1 \myidu/_1676_ ( .D(\myidu/_0946_ ), .CK(clock ), .Q(\ID_EX_typ [6] ), .QN(\myidu/_0865_ ) );
DFF_X1 \myidu/_1677_ ( .D(\myidu/_0947_ ), .CK(clock ), .Q(\ID_EX_typ [7] ), .QN(\myidu/_0864_ ) );
DFF_X1 \myidu/_1678_ ( .D(\myidu/_0948_ ), .CK(clock ), .Q(\ID_EX_pc [0] ), .QN(\myidu/_0863_ ) );
DFF_X1 \myidu/_1679_ ( .D(\myidu/_0949_ ), .CK(clock ), .Q(\ID_EX_pc [1] ), .QN(\myidu/_0862_ ) );
DFF_X1 \myidu/_1680_ ( .D(\myidu/_0950_ ), .CK(clock ), .Q(\ID_EX_pc [2] ), .QN(\myidu/_0861_ ) );
DFF_X1 \myidu/_1681_ ( .D(\myidu/_0951_ ), .CK(clock ), .Q(\ID_EX_pc [3] ), .QN(\myidu/_0860_ ) );
DFF_X1 \myidu/_1682_ ( .D(\myidu/_0952_ ), .CK(clock ), .Q(\ID_EX_pc [4] ), .QN(\myidu/_0859_ ) );
DFF_X1 \myidu/_1683_ ( .D(\myidu/_0953_ ), .CK(clock ), .Q(\ID_EX_pc [5] ), .QN(\myidu/_0858_ ) );
DFF_X1 \myidu/_1684_ ( .D(\myidu/_0954_ ), .CK(clock ), .Q(\ID_EX_pc [6] ), .QN(\myidu/_0857_ ) );
DFF_X1 \myidu/_1685_ ( .D(\myidu/_0955_ ), .CK(clock ), .Q(\ID_EX_pc [7] ), .QN(\myidu/_0856_ ) );
DFF_X1 \myidu/_1686_ ( .D(\myidu/_0956_ ), .CK(clock ), .Q(\ID_EX_pc [8] ), .QN(\myidu/_0855_ ) );
DFF_X1 \myidu/_1687_ ( .D(\myidu/_0957_ ), .CK(clock ), .Q(\ID_EX_pc [9] ), .QN(\myidu/_0854_ ) );
DFF_X1 \myidu/_1688_ ( .D(\myidu/_0958_ ), .CK(clock ), .Q(\ID_EX_pc [10] ), .QN(\myidu/_0853_ ) );
DFF_X1 \myidu/_1689_ ( .D(\myidu/_0959_ ), .CK(clock ), .Q(\ID_EX_pc [11] ), .QN(\myidu/_0852_ ) );
DFF_X1 \myidu/_1690_ ( .D(\myidu/_0960_ ), .CK(clock ), .Q(\ID_EX_pc [12] ), .QN(\myidu/_0851_ ) );
DFF_X1 \myidu/_1691_ ( .D(\myidu/_0961_ ), .CK(clock ), .Q(\ID_EX_pc [13] ), .QN(\myidu/_0850_ ) );
DFF_X1 \myidu/_1692_ ( .D(\myidu/_0962_ ), .CK(clock ), .Q(\ID_EX_pc [14] ), .QN(\myidu/_0849_ ) );
DFF_X1 \myidu/_1693_ ( .D(\myidu/_0963_ ), .CK(clock ), .Q(\ID_EX_pc [15] ), .QN(\myidu/_0848_ ) );
DFF_X1 \myidu/_1694_ ( .D(\myidu/_0964_ ), .CK(clock ), .Q(\ID_EX_pc [16] ), .QN(\myidu/_0847_ ) );
DFF_X1 \myidu/_1695_ ( .D(\myidu/_0965_ ), .CK(clock ), .Q(\ID_EX_pc [17] ), .QN(\myidu/_0846_ ) );
DFF_X1 \myidu/_1696_ ( .D(\myidu/_0966_ ), .CK(clock ), .Q(\ID_EX_pc [18] ), .QN(\myidu/_0845_ ) );
DFF_X1 \myidu/_1697_ ( .D(\myidu/_0967_ ), .CK(clock ), .Q(\ID_EX_pc [19] ), .QN(\myidu/_0844_ ) );
DFF_X1 \myidu/_1698_ ( .D(\myidu/_0968_ ), .CK(clock ), .Q(\ID_EX_pc [20] ), .QN(\myidu/_0843_ ) );
DFF_X1 \myidu/_1699_ ( .D(\myidu/_0969_ ), .CK(clock ), .Q(\ID_EX_pc [21] ), .QN(\myidu/_0842_ ) );
DFF_X1 \myidu/_1700_ ( .D(\myidu/_0970_ ), .CK(clock ), .Q(\ID_EX_pc [22] ), .QN(\myidu/_0841_ ) );
DFF_X1 \myidu/_1701_ ( .D(\myidu/_0971_ ), .CK(clock ), .Q(\ID_EX_pc [23] ), .QN(\myidu/_0840_ ) );
DFF_X1 \myidu/_1702_ ( .D(\myidu/_0972_ ), .CK(clock ), .Q(\ID_EX_pc [24] ), .QN(\myidu/_0839_ ) );
DFF_X1 \myidu/_1703_ ( .D(\myidu/_0973_ ), .CK(clock ), .Q(\ID_EX_pc [25] ), .QN(\myidu/_0838_ ) );
DFF_X1 \myidu/_1704_ ( .D(\myidu/_0974_ ), .CK(clock ), .Q(\ID_EX_pc [26] ), .QN(\myidu/_0837_ ) );
DFF_X1 \myidu/_1705_ ( .D(\myidu/_0975_ ), .CK(clock ), .Q(\ID_EX_pc [27] ), .QN(\myidu/_0836_ ) );
DFF_X1 \myidu/_1706_ ( .D(\myidu/_0976_ ), .CK(clock ), .Q(\ID_EX_pc [28] ), .QN(\myidu/_0835_ ) );
DFF_X1 \myidu/_1707_ ( .D(\myidu/_0977_ ), .CK(clock ), .Q(\ID_EX_pc [29] ), .QN(\myidu/_0834_ ) );
DFF_X1 \myidu/_1708_ ( .D(\myidu/_0978_ ), .CK(clock ), .Q(\ID_EX_pc [30] ), .QN(\myidu/_0833_ ) );
DFF_X1 \myidu/_1709_ ( .D(\myidu/_0979_ ), .CK(clock ), .Q(\ID_EX_pc [31] ), .QN(\myidu/_0832_ ) );
DFF_X1 \myidu/_1710_ ( .D(\myidu/_0980_ ), .CK(clock ), .Q(\ID_EX_rs1 [0] ), .QN(\myidu/_0831_ ) );
DFF_X1 \myidu/_1711_ ( .D(\myidu/_0981_ ), .CK(clock ), .Q(\ID_EX_rs1 [1] ), .QN(\myidu/_0830_ ) );
DFF_X1 \myidu/_1712_ ( .D(\myidu/_0982_ ), .CK(clock ), .Q(\ID_EX_rs1 [2] ), .QN(\myidu/_0829_ ) );
DFF_X1 \myidu/_1713_ ( .D(\myidu/_0983_ ), .CK(clock ), .Q(\ID_EX_rs1 [3] ), .QN(\myidu/_0828_ ) );
DFF_X1 \myidu/_1714_ ( .D(\myidu/_0984_ ), .CK(clock ), .Q(\ID_EX_rs1 [4] ), .QN(\myidu/_0827_ ) );
DFF_X1 \myidu/_1715_ ( .D(\myidu/_0985_ ), .CK(clock ), .Q(\ID_EX_rs2 [0] ), .QN(\myidu/_0826_ ) );
DFF_X1 \myidu/_1716_ ( .D(\myidu/_0986_ ), .CK(clock ), .Q(\ID_EX_rs2 [1] ), .QN(\myidu/_0825_ ) );
DFF_X1 \myidu/_1717_ ( .D(\myidu/_0987_ ), .CK(clock ), .Q(\ID_EX_rs2 [2] ), .QN(\myidu/_0824_ ) );
DFF_X1 \myidu/_1718_ ( .D(\myidu/_0988_ ), .CK(clock ), .Q(\ID_EX_rs2 [3] ), .QN(\myidu/_0823_ ) );
DFF_X1 \myidu/_1719_ ( .D(\myidu/_0989_ ), .CK(clock ), .Q(\ID_EX_rs2 [4] ), .QN(\myidu/_0822_ ) );
DFF_X1 \myidu/_1720_ ( .D(\myidu/_0990_ ), .CK(clock ), .Q(\ID_EX_rd [0] ), .QN(\myidu/_0821_ ) );
DFF_X1 \myidu/_1721_ ( .D(\myidu/_0991_ ), .CK(clock ), .Q(\ID_EX_rd [1] ), .QN(\myidu/_0820_ ) );
DFF_X1 \myidu/_1722_ ( .D(\myidu/_0992_ ), .CK(clock ), .Q(\ID_EX_rd [2] ), .QN(\myidu/_0819_ ) );
DFF_X1 \myidu/_1723_ ( .D(\myidu/_0993_ ), .CK(clock ), .Q(\ID_EX_rd [3] ), .QN(\myidu/_0818_ ) );
DFF_X1 \myidu/_1724_ ( .D(\myidu/_0994_ ), .CK(clock ), .Q(\ID_EX_rd [4] ), .QN(\myidu/_0817_ ) );
DFF_X1 \myidu/_1725_ ( .D(\myidu/_0995_ ), .CK(clock ), .Q(\ID_EX_csr [0] ), .QN(\myidu/_0816_ ) );
DFF_X1 \myidu/_1726_ ( .D(\myidu/_0996_ ), .CK(clock ), .Q(\ID_EX_csr [1] ), .QN(\myidu/_0815_ ) );
DFF_X1 \myidu/_1727_ ( .D(\myidu/_0997_ ), .CK(clock ), .Q(\ID_EX_csr [2] ), .QN(\myidu/_0814_ ) );
DFF_X1 \myidu/_1728_ ( .D(\myidu/_0998_ ), .CK(clock ), .Q(\ID_EX_csr [3] ), .QN(\myidu/_0813_ ) );
DFF_X1 \myidu/_1729_ ( .D(\myidu/_0999_ ), .CK(clock ), .Q(\ID_EX_csr [4] ), .QN(\myidu/_0812_ ) );
DFF_X1 \myidu/_1730_ ( .D(\myidu/_1000_ ), .CK(clock ), .Q(\ID_EX_csr [5] ), .QN(\myidu/_0811_ ) );
DFF_X1 \myidu/_1731_ ( .D(\myidu/_1001_ ), .CK(clock ), .Q(\ID_EX_csr [6] ), .QN(\myidu/_0810_ ) );
DFF_X1 \myidu/_1732_ ( .D(\myidu/_1002_ ), .CK(clock ), .Q(\ID_EX_csr [7] ), .QN(\myidu/_0809_ ) );
DFF_X1 \myidu/_1733_ ( .D(\myidu/_1003_ ), .CK(clock ), .Q(\ID_EX_csr [8] ), .QN(\myidu/_0808_ ) );
DFF_X1 \myidu/_1734_ ( .D(\myidu/_1004_ ), .CK(clock ), .Q(\ID_EX_csr [9] ), .QN(\myidu/_0807_ ) );
DFF_X1 \myidu/_1735_ ( .D(\myidu/_1005_ ), .CK(clock ), .Q(\ID_EX_csr [10] ), .QN(\myidu/_0806_ ) );
DFF_X1 \myidu/_1736_ ( .D(\myidu/_1006_ ), .CK(clock ), .Q(\ID_EX_csr [11] ), .QN(\myidu/_0805_ ) );
DFF_X1 \myidu/_1737_ ( .D(\myidu/_1007_ ), .CK(clock ), .Q(stall_quest_loaduse ), .QN(\myidu/_0804_ ) );
DFF_X1 \myidu/_1738_ ( .D(\myidu/_1008_ ), .CK(clock ), .Q(fc_disenable ), .QN(\myidu/_0803_ ) );
BUF_X1 \myidu/_1739_ ( .A(IDU_ready_IFU ), .Z(\myidu/state [0] ) );
BUF_X1 \myidu/_1740_ ( .A(IDU_valid_EXU ), .Z(\myidu/state [1] ) );
BUF_X1 \myidu/_1741_ ( .A(\ID_EX_typ [6] ), .Z(\myidu/_0799_ ) );
BUF_X1 \myidu/_1742_ ( .A(\ID_EX_typ [5] ), .Z(\myidu/_0798_ ) );
BUF_X1 \myidu/_1743_ ( .A(\ID_EX_typ [7] ), .Z(\myidu/_0800_ ) );
BUF_X1 \myidu/_1744_ ( .A(\IF_ID_inst [15] ), .Z(\myidu/_0161_ ) );
BUF_X1 \myidu/_1745_ ( .A(\ID_EX_rd [0] ), .Z(\myidu/_0772_ ) );
BUF_X1 \myidu/_1746_ ( .A(\IF_ID_inst [16] ), .Z(\myidu/_0162_ ) );
BUF_X1 \myidu/_1747_ ( .A(\ID_EX_rd [1] ), .Z(\myidu/_0773_ ) );
BUF_X1 \myidu/_1748_ ( .A(\IF_ID_inst [17] ), .Z(\myidu/_0163_ ) );
BUF_X1 \myidu/_1749_ ( .A(\ID_EX_rd [2] ), .Z(\myidu/_0774_ ) );
BUF_X1 \myidu/_1750_ ( .A(\IF_ID_inst [18] ), .Z(\myidu/_0164_ ) );
BUF_X1 \myidu/_1751_ ( .A(\ID_EX_rd [3] ), .Z(\myidu/_0775_ ) );
BUF_X1 \myidu/_1752_ ( .A(\IF_ID_inst [19] ), .Z(\myidu/_0165_ ) );
BUF_X1 \myidu/_1753_ ( .A(\ID_EX_rd [4] ), .Z(\myidu/_0776_ ) );
BUF_X1 \myidu/_1754_ ( .A(\IF_ID_inst [20] ), .Z(\myidu/_0167_ ) );
BUF_X1 \myidu/_1755_ ( .A(\IF_ID_inst [21] ), .Z(\myidu/_0168_ ) );
BUF_X1 \myidu/_1756_ ( .A(\IF_ID_inst [22] ), .Z(\myidu/_0169_ ) );
BUF_X1 \myidu/_1757_ ( .A(\IF_ID_inst [23] ), .Z(\myidu/_0170_ ) );
BUF_X1 \myidu/_1758_ ( .A(\IF_ID_inst [24] ), .Z(\myidu/_0171_ ) );
BUF_X1 \myidu/_1759_ ( .A(\IF_ID_inst [1] ), .Z(\myidu/_0166_ ) );
BUF_X1 \myidu/_1760_ ( .A(\IF_ID_inst [0] ), .Z(\myidu/_0155_ ) );
BUF_X1 \myidu/_1761_ ( .A(\IF_ID_inst [3] ), .Z(\myidu/_0180_ ) );
BUF_X1 \myidu/_1762_ ( .A(\IF_ID_inst [2] ), .Z(\myidu/_0177_ ) );
BUF_X1 \myidu/_1763_ ( .A(\IF_ID_inst [5] ), .Z(\myidu/_0182_ ) );
BUF_X1 \myidu/_1764_ ( .A(\IF_ID_inst [4] ), .Z(\myidu/_0181_ ) );
BUF_X1 \myidu/_1765_ ( .A(\IF_ID_inst [6] ), .Z(\myidu/_0183_ ) );
BUF_X1 \myidu/_1766_ ( .A(\IF_ID_inst [12] ), .Z(\myidu/_0158_ ) );
BUF_X1 \myidu/_1767_ ( .A(\IF_ID_inst [14] ), .Z(\myidu/_0160_ ) );
BUF_X1 \myidu/_1768_ ( .A(\IF_ID_inst [13] ), .Z(\myidu/_0159_ ) );
BUF_X1 \myidu/_1769_ ( .A(\IF_ID_inst [7] ), .Z(\myidu/_0184_ ) );
BUF_X1 \myidu/_1770_ ( .A(\IF_ID_inst [9] ), .Z(\myidu/_0186_ ) );
BUF_X1 \myidu/_1771_ ( .A(\IF_ID_inst [8] ), .Z(\myidu/_0185_ ) );
BUF_X1 \myidu/_1772_ ( .A(\IF_ID_inst [11] ), .Z(\myidu/_0157_ ) );
BUF_X1 \myidu/_1773_ ( .A(\IF_ID_inst [10] ), .Z(\myidu/_0156_ ) );
BUF_X1 \myidu/_1774_ ( .A(\IF_ID_inst [25] ), .Z(\myidu/_0172_ ) );
BUF_X1 \myidu/_1775_ ( .A(\IF_ID_inst [27] ), .Z(\myidu/_0174_ ) );
BUF_X1 \myidu/_1776_ ( .A(\IF_ID_inst [26] ), .Z(\myidu/_0173_ ) );
BUF_X1 \myidu/_1777_ ( .A(\IF_ID_inst [29] ), .Z(\myidu/_0176_ ) );
BUF_X1 \myidu/_1778_ ( .A(\IF_ID_inst [28] ), .Z(\myidu/_0175_ ) );
BUF_X1 \myidu/_1779_ ( .A(\IF_ID_inst [31] ), .Z(\myidu/_0179_ ) );
BUF_X1 \myidu/_1780_ ( .A(\IF_ID_inst [30] ), .Z(\myidu/_0178_ ) );
BUF_X1 \myidu/_1781_ ( .A(IDU_ready_IFU ), .Z(\myidu/_0778_ ) );
BUF_X1 \myidu/_1782_ ( .A(reset ), .Z(\myidu/_0789_ ) );
BUF_X1 \myidu/_1783_ ( .A(IFU_valid_IDU ), .Z(\myidu/_0801_ ) );
BUF_X1 \myidu/_1784_ ( .A(EXU_ready_IDU ), .Z(\myidu/_0777_ ) );
BUF_X1 \myidu/_1785_ ( .A(IDU_valid_EXU ), .Z(\myidu/_0802_ ) );
BUF_X1 \myidu/_1786_ ( .A(loaduse_clear ), .Z(\myidu/_0187_ ) );
BUF_X1 \myidu/_1787_ ( .A(\myidu/state [2] ), .Z(\myidu/_0792_ ) );
BUF_X1 \myidu/_1788_ ( .A(\myidu/_0005_ ), .Z(\myidu/_0001_ ) );
BUF_X1 \myidu/_1789_ ( .A(\myidu/_0004_ ), .Z(\myidu/_0000_ ) );
BUF_X1 \myidu/_1790_ ( .A(\myidu/_0006_ ), .Z(\myidu/_0002_ ) );
BUF_X1 \myidu/_1791_ ( .A(\myidu/_0003_ ), .Z(\myidu/_0007_ ) );
BUF_X1 \myidu/_1792_ ( .A(\ID_EX_imm [0] ), .Z(\myidu/_0123_ ) );
BUF_X1 \myidu/_1793_ ( .A(\myidu/_0008_ ), .Z(\myidu/_0907_ ) );
BUF_X1 \myidu/_1794_ ( .A(\ID_EX_imm [1] ), .Z(\myidu/_0134_ ) );
BUF_X1 \myidu/_1795_ ( .A(\myidu/_0009_ ), .Z(\myidu/_0908_ ) );
BUF_X1 \myidu/_1796_ ( .A(\ID_EX_imm [2] ), .Z(\myidu/_0145_ ) );
BUF_X1 \myidu/_1797_ ( .A(\myidu/_0010_ ), .Z(\myidu/_0909_ ) );
BUF_X1 \myidu/_1798_ ( .A(\ID_EX_imm [3] ), .Z(\myidu/_0148_ ) );
BUF_X1 \myidu/_1799_ ( .A(\myidu/_0011_ ), .Z(\myidu/_0910_ ) );
BUF_X1 \myidu/_1800_ ( .A(\ID_EX_imm [4] ), .Z(\myidu/_0149_ ) );
BUF_X1 \myidu/_1801_ ( .A(\myidu/_0012_ ), .Z(\myidu/_0911_ ) );
BUF_X1 \myidu/_1802_ ( .A(\ID_EX_imm [5] ), .Z(\myidu/_0150_ ) );
BUF_X1 \myidu/_1803_ ( .A(\myidu/_0013_ ), .Z(\myidu/_0912_ ) );
BUF_X1 \myidu/_1804_ ( .A(\ID_EX_imm [6] ), .Z(\myidu/_0151_ ) );
BUF_X1 \myidu/_1805_ ( .A(\myidu/_0014_ ), .Z(\myidu/_0913_ ) );
BUF_X1 \myidu/_1806_ ( .A(\ID_EX_imm [7] ), .Z(\myidu/_0152_ ) );
BUF_X1 \myidu/_1807_ ( .A(\myidu/_0015_ ), .Z(\myidu/_0914_ ) );
BUF_X1 \myidu/_1808_ ( .A(\ID_EX_imm [8] ), .Z(\myidu/_0153_ ) );
BUF_X1 \myidu/_1809_ ( .A(\myidu/_0016_ ), .Z(\myidu/_0915_ ) );
BUF_X1 \myidu/_1810_ ( .A(\ID_EX_imm [9] ), .Z(\myidu/_0154_ ) );
BUF_X1 \myidu/_1811_ ( .A(\myidu/_0017_ ), .Z(\myidu/_0916_ ) );
BUF_X1 \myidu/_1812_ ( .A(\ID_EX_imm [10] ), .Z(\myidu/_0124_ ) );
BUF_X1 \myidu/_1813_ ( .A(\myidu/_0018_ ), .Z(\myidu/_0917_ ) );
BUF_X1 \myidu/_1814_ ( .A(\ID_EX_imm [11] ), .Z(\myidu/_0125_ ) );
BUF_X1 \myidu/_1815_ ( .A(\myidu/_0019_ ), .Z(\myidu/_0918_ ) );
BUF_X1 \myidu/_1816_ ( .A(\ID_EX_imm [12] ), .Z(\myidu/_0126_ ) );
BUF_X1 \myidu/_1817_ ( .A(\myidu/_0020_ ), .Z(\myidu/_0919_ ) );
BUF_X1 \myidu/_1818_ ( .A(\ID_EX_imm [13] ), .Z(\myidu/_0127_ ) );
BUF_X1 \myidu/_1819_ ( .A(\myidu/_0021_ ), .Z(\myidu/_0920_ ) );
BUF_X1 \myidu/_1820_ ( .A(\ID_EX_imm [14] ), .Z(\myidu/_0128_ ) );
BUF_X1 \myidu/_1821_ ( .A(\myidu/_0022_ ), .Z(\myidu/_0921_ ) );
BUF_X1 \myidu/_1822_ ( .A(\ID_EX_imm [15] ), .Z(\myidu/_0129_ ) );
BUF_X1 \myidu/_1823_ ( .A(\myidu/_0023_ ), .Z(\myidu/_0922_ ) );
BUF_X1 \myidu/_1824_ ( .A(\ID_EX_imm [16] ), .Z(\myidu/_0130_ ) );
BUF_X1 \myidu/_1825_ ( .A(\myidu/_0024_ ), .Z(\myidu/_0923_ ) );
BUF_X1 \myidu/_1826_ ( .A(\ID_EX_imm [17] ), .Z(\myidu/_0131_ ) );
BUF_X1 \myidu/_1827_ ( .A(\myidu/_0025_ ), .Z(\myidu/_0924_ ) );
BUF_X1 \myidu/_1828_ ( .A(\ID_EX_imm [18] ), .Z(\myidu/_0132_ ) );
BUF_X1 \myidu/_1829_ ( .A(\myidu/_0026_ ), .Z(\myidu/_0925_ ) );
BUF_X1 \myidu/_1830_ ( .A(\ID_EX_imm [19] ), .Z(\myidu/_0133_ ) );
BUF_X1 \myidu/_1831_ ( .A(\myidu/_0027_ ), .Z(\myidu/_0926_ ) );
BUF_X1 \myidu/_1832_ ( .A(\ID_EX_imm [20] ), .Z(\myidu/_0135_ ) );
BUF_X1 \myidu/_1833_ ( .A(\myidu/_0028_ ), .Z(\myidu/_0927_ ) );
BUF_X1 \myidu/_1834_ ( .A(\ID_EX_imm [21] ), .Z(\myidu/_0136_ ) );
BUF_X1 \myidu/_1835_ ( .A(\myidu/_0029_ ), .Z(\myidu/_0928_ ) );
BUF_X1 \myidu/_1836_ ( .A(\ID_EX_imm [22] ), .Z(\myidu/_0137_ ) );
BUF_X1 \myidu/_1837_ ( .A(\myidu/_0030_ ), .Z(\myidu/_0929_ ) );
BUF_X1 \myidu/_1838_ ( .A(\ID_EX_imm [23] ), .Z(\myidu/_0138_ ) );
BUF_X1 \myidu/_1839_ ( .A(\myidu/_0031_ ), .Z(\myidu/_0930_ ) );
BUF_X1 \myidu/_1840_ ( .A(\ID_EX_imm [24] ), .Z(\myidu/_0139_ ) );
BUF_X1 \myidu/_1841_ ( .A(\myidu/_0032_ ), .Z(\myidu/_0931_ ) );
BUF_X1 \myidu/_1842_ ( .A(\ID_EX_imm [25] ), .Z(\myidu/_0140_ ) );
BUF_X1 \myidu/_1843_ ( .A(\myidu/_0033_ ), .Z(\myidu/_0932_ ) );
BUF_X1 \myidu/_1844_ ( .A(\ID_EX_imm [26] ), .Z(\myidu/_0141_ ) );
BUF_X1 \myidu/_1845_ ( .A(\myidu/_0034_ ), .Z(\myidu/_0933_ ) );
BUF_X1 \myidu/_1846_ ( .A(\ID_EX_imm [27] ), .Z(\myidu/_0142_ ) );
BUF_X1 \myidu/_1847_ ( .A(\myidu/_0035_ ), .Z(\myidu/_0934_ ) );
BUF_X1 \myidu/_1848_ ( .A(\ID_EX_imm [28] ), .Z(\myidu/_0143_ ) );
BUF_X1 \myidu/_1849_ ( .A(\myidu/_0036_ ), .Z(\myidu/_0935_ ) );
BUF_X1 \myidu/_1850_ ( .A(\ID_EX_imm [29] ), .Z(\myidu/_0144_ ) );
BUF_X1 \myidu/_1851_ ( .A(\myidu/_0037_ ), .Z(\myidu/_0936_ ) );
BUF_X1 \myidu/_1852_ ( .A(\ID_EX_imm [30] ), .Z(\myidu/_0146_ ) );
BUF_X1 \myidu/_1853_ ( .A(\myidu/_0038_ ), .Z(\myidu/_0937_ ) );
BUF_X1 \myidu/_1854_ ( .A(\ID_EX_imm [31] ), .Z(\myidu/_0147_ ) );
BUF_X1 \myidu/_1855_ ( .A(\myidu/_0039_ ), .Z(\myidu/_0938_ ) );
BUF_X1 \myidu/_1856_ ( .A(stall_quest_fencei ), .Z(\myidu/_0790_ ) );
BUF_X1 \myidu/_1857_ ( .A(\ID_EX_typ [0] ), .Z(\myidu/_0793_ ) );
BUF_X1 \myidu/_1858_ ( .A(\ID_EX_typ [1] ), .Z(\myidu/_0794_ ) );
BUF_X1 \myidu/_1859_ ( .A(\ID_EX_typ [2] ), .Z(\myidu/_0795_ ) );
BUF_X1 \myidu/_1860_ ( .A(\ID_EX_typ [3] ), .Z(\myidu/_0796_ ) );
BUF_X1 \myidu/_1861_ ( .A(\ID_EX_typ [4] ), .Z(\myidu/_0797_ ) );
BUF_X1 \myidu/_1862_ ( .A(\ID_EX_pc [0] ), .Z(\myidu/_0740_ ) );
BUF_X1 \myidu/_1863_ ( .A(\IF_ID_pc [0] ), .Z(\myidu/_0708_ ) );
BUF_X1 \myidu/_1864_ ( .A(\myidu/_0049_ ), .Z(\myidu/_0948_ ) );
BUF_X1 \myidu/_1865_ ( .A(\ID_EX_pc [1] ), .Z(\myidu/_0751_ ) );
BUF_X1 \myidu/_1866_ ( .A(\IF_ID_pc [1] ), .Z(\myidu/_0719_ ) );
BUF_X1 \myidu/_1867_ ( .A(\myidu/_0050_ ), .Z(\myidu/_0949_ ) );
BUF_X1 \myidu/_1868_ ( .A(\ID_EX_pc [2] ), .Z(\myidu/_0762_ ) );
BUF_X1 \myidu/_1869_ ( .A(\IF_ID_pc [2] ), .Z(\myidu/_0730_ ) );
BUF_X1 \myidu/_1870_ ( .A(\myidu/_0051_ ), .Z(\myidu/_0950_ ) );
BUF_X1 \myidu/_1871_ ( .A(\ID_EX_pc [3] ), .Z(\myidu/_0765_ ) );
BUF_X1 \myidu/_1872_ ( .A(\IF_ID_pc [3] ), .Z(\myidu/_0733_ ) );
BUF_X1 \myidu/_1873_ ( .A(\myidu/_0052_ ), .Z(\myidu/_0951_ ) );
BUF_X1 \myidu/_1874_ ( .A(\ID_EX_pc [4] ), .Z(\myidu/_0766_ ) );
BUF_X1 \myidu/_1875_ ( .A(\IF_ID_pc [4] ), .Z(\myidu/_0734_ ) );
BUF_X1 \myidu/_1876_ ( .A(\myidu/_0053_ ), .Z(\myidu/_0952_ ) );
BUF_X1 \myidu/_1877_ ( .A(\ID_EX_pc [5] ), .Z(\myidu/_0767_ ) );
BUF_X1 \myidu/_1878_ ( .A(\IF_ID_pc [5] ), .Z(\myidu/_0735_ ) );
BUF_X1 \myidu/_1879_ ( .A(\myidu/_0054_ ), .Z(\myidu/_0953_ ) );
BUF_X1 \myidu/_1880_ ( .A(\ID_EX_pc [6] ), .Z(\myidu/_0768_ ) );
BUF_X1 \myidu/_1881_ ( .A(\IF_ID_pc [6] ), .Z(\myidu/_0736_ ) );
BUF_X1 \myidu/_1882_ ( .A(\myidu/_0055_ ), .Z(\myidu/_0954_ ) );
BUF_X1 \myidu/_1883_ ( .A(\ID_EX_pc [7] ), .Z(\myidu/_0769_ ) );
BUF_X1 \myidu/_1884_ ( .A(\IF_ID_pc [7] ), .Z(\myidu/_0737_ ) );
BUF_X1 \myidu/_1885_ ( .A(\myidu/_0056_ ), .Z(\myidu/_0955_ ) );
BUF_X1 \myidu/_1886_ ( .A(\ID_EX_pc [8] ), .Z(\myidu/_0770_ ) );
BUF_X1 \myidu/_1887_ ( .A(\IF_ID_pc [8] ), .Z(\myidu/_0738_ ) );
BUF_X1 \myidu/_1888_ ( .A(\myidu/_0057_ ), .Z(\myidu/_0956_ ) );
BUF_X1 \myidu/_1889_ ( .A(\ID_EX_pc [9] ), .Z(\myidu/_0771_ ) );
BUF_X1 \myidu/_1890_ ( .A(\IF_ID_pc [9] ), .Z(\myidu/_0739_ ) );
BUF_X1 \myidu/_1891_ ( .A(\myidu/_0058_ ), .Z(\myidu/_0957_ ) );
BUF_X1 \myidu/_1892_ ( .A(\ID_EX_pc [10] ), .Z(\myidu/_0741_ ) );
BUF_X1 \myidu/_1893_ ( .A(\IF_ID_pc [10] ), .Z(\myidu/_0709_ ) );
BUF_X1 \myidu/_1894_ ( .A(\myidu/_0059_ ), .Z(\myidu/_0958_ ) );
BUF_X1 \myidu/_1895_ ( .A(\ID_EX_pc [11] ), .Z(\myidu/_0742_ ) );
BUF_X1 \myidu/_1896_ ( .A(\IF_ID_pc [11] ), .Z(\myidu/_0710_ ) );
BUF_X1 \myidu/_1897_ ( .A(\myidu/_0060_ ), .Z(\myidu/_0959_ ) );
BUF_X1 \myidu/_1898_ ( .A(\ID_EX_pc [12] ), .Z(\myidu/_0743_ ) );
BUF_X1 \myidu/_1899_ ( .A(\IF_ID_pc [12] ), .Z(\myidu/_0711_ ) );
BUF_X1 \myidu/_1900_ ( .A(\myidu/_0061_ ), .Z(\myidu/_0960_ ) );
BUF_X1 \myidu/_1901_ ( .A(\ID_EX_pc [13] ), .Z(\myidu/_0744_ ) );
BUF_X1 \myidu/_1902_ ( .A(\IF_ID_pc [13] ), .Z(\myidu/_0712_ ) );
BUF_X1 \myidu/_1903_ ( .A(\myidu/_0062_ ), .Z(\myidu/_0961_ ) );
BUF_X1 \myidu/_1904_ ( .A(\ID_EX_pc [14] ), .Z(\myidu/_0745_ ) );
BUF_X1 \myidu/_1905_ ( .A(\IF_ID_pc [14] ), .Z(\myidu/_0713_ ) );
BUF_X1 \myidu/_1906_ ( .A(\myidu/_0063_ ), .Z(\myidu/_0962_ ) );
BUF_X1 \myidu/_1907_ ( .A(\ID_EX_pc [15] ), .Z(\myidu/_0746_ ) );
BUF_X1 \myidu/_1908_ ( .A(\IF_ID_pc [15] ), .Z(\myidu/_0714_ ) );
BUF_X1 \myidu/_1909_ ( .A(\myidu/_0064_ ), .Z(\myidu/_0963_ ) );
BUF_X1 \myidu/_1910_ ( .A(\ID_EX_pc [16] ), .Z(\myidu/_0747_ ) );
BUF_X1 \myidu/_1911_ ( .A(\IF_ID_pc [16] ), .Z(\myidu/_0715_ ) );
BUF_X1 \myidu/_1912_ ( .A(\myidu/_0065_ ), .Z(\myidu/_0964_ ) );
BUF_X1 \myidu/_1913_ ( .A(\ID_EX_pc [17] ), .Z(\myidu/_0748_ ) );
BUF_X1 \myidu/_1914_ ( .A(\IF_ID_pc [17] ), .Z(\myidu/_0716_ ) );
BUF_X1 \myidu/_1915_ ( .A(\myidu/_0066_ ), .Z(\myidu/_0965_ ) );
BUF_X1 \myidu/_1916_ ( .A(\ID_EX_pc [18] ), .Z(\myidu/_0749_ ) );
BUF_X1 \myidu/_1917_ ( .A(\IF_ID_pc [18] ), .Z(\myidu/_0717_ ) );
BUF_X1 \myidu/_1918_ ( .A(\myidu/_0067_ ), .Z(\myidu/_0966_ ) );
BUF_X1 \myidu/_1919_ ( .A(\ID_EX_pc [19] ), .Z(\myidu/_0750_ ) );
BUF_X1 \myidu/_1920_ ( .A(\IF_ID_pc [19] ), .Z(\myidu/_0718_ ) );
BUF_X1 \myidu/_1921_ ( .A(\myidu/_0068_ ), .Z(\myidu/_0967_ ) );
BUF_X1 \myidu/_1922_ ( .A(\ID_EX_pc [20] ), .Z(\myidu/_0752_ ) );
BUF_X1 \myidu/_1923_ ( .A(\IF_ID_pc [20] ), .Z(\myidu/_0720_ ) );
BUF_X1 \myidu/_1924_ ( .A(\myidu/_0069_ ), .Z(\myidu/_0968_ ) );
BUF_X1 \myidu/_1925_ ( .A(\ID_EX_pc [21] ), .Z(\myidu/_0753_ ) );
BUF_X1 \myidu/_1926_ ( .A(\IF_ID_pc [21] ), .Z(\myidu/_0721_ ) );
BUF_X1 \myidu/_1927_ ( .A(\myidu/_0070_ ), .Z(\myidu/_0969_ ) );
BUF_X1 \myidu/_1928_ ( .A(\ID_EX_pc [22] ), .Z(\myidu/_0754_ ) );
BUF_X1 \myidu/_1929_ ( .A(\IF_ID_pc [22] ), .Z(\myidu/_0722_ ) );
BUF_X1 \myidu/_1930_ ( .A(\myidu/_0071_ ), .Z(\myidu/_0970_ ) );
BUF_X1 \myidu/_1931_ ( .A(\ID_EX_pc [23] ), .Z(\myidu/_0755_ ) );
BUF_X1 \myidu/_1932_ ( .A(\IF_ID_pc [23] ), .Z(\myidu/_0723_ ) );
BUF_X1 \myidu/_1933_ ( .A(\myidu/_0072_ ), .Z(\myidu/_0971_ ) );
BUF_X1 \myidu/_1934_ ( .A(\ID_EX_pc [24] ), .Z(\myidu/_0756_ ) );
BUF_X1 \myidu/_1935_ ( .A(\IF_ID_pc [24] ), .Z(\myidu/_0724_ ) );
BUF_X1 \myidu/_1936_ ( .A(\myidu/_0073_ ), .Z(\myidu/_0972_ ) );
BUF_X1 \myidu/_1937_ ( .A(\ID_EX_pc [25] ), .Z(\myidu/_0757_ ) );
BUF_X1 \myidu/_1938_ ( .A(\IF_ID_pc [25] ), .Z(\myidu/_0725_ ) );
BUF_X1 \myidu/_1939_ ( .A(\myidu/_0074_ ), .Z(\myidu/_0973_ ) );
BUF_X1 \myidu/_1940_ ( .A(\ID_EX_pc [26] ), .Z(\myidu/_0758_ ) );
BUF_X1 \myidu/_1941_ ( .A(\IF_ID_pc [26] ), .Z(\myidu/_0726_ ) );
BUF_X1 \myidu/_1942_ ( .A(\myidu/_0075_ ), .Z(\myidu/_0974_ ) );
BUF_X1 \myidu/_1943_ ( .A(\ID_EX_pc [27] ), .Z(\myidu/_0759_ ) );
BUF_X1 \myidu/_1944_ ( .A(\IF_ID_pc [27] ), .Z(\myidu/_0727_ ) );
BUF_X1 \myidu/_1945_ ( .A(\myidu/_0076_ ), .Z(\myidu/_0975_ ) );
BUF_X1 \myidu/_1946_ ( .A(\ID_EX_pc [28] ), .Z(\myidu/_0760_ ) );
BUF_X1 \myidu/_1947_ ( .A(\IF_ID_pc [28] ), .Z(\myidu/_0728_ ) );
BUF_X1 \myidu/_1948_ ( .A(\myidu/_0077_ ), .Z(\myidu/_0976_ ) );
BUF_X1 \myidu/_1949_ ( .A(\ID_EX_pc [29] ), .Z(\myidu/_0761_ ) );
BUF_X1 \myidu/_1950_ ( .A(\IF_ID_pc [29] ), .Z(\myidu/_0729_ ) );
BUF_X1 \myidu/_1951_ ( .A(\myidu/_0078_ ), .Z(\myidu/_0977_ ) );
BUF_X1 \myidu/_1952_ ( .A(\ID_EX_pc [30] ), .Z(\myidu/_0763_ ) );
BUF_X1 \myidu/_1953_ ( .A(\IF_ID_pc [30] ), .Z(\myidu/_0731_ ) );
BUF_X1 \myidu/_1954_ ( .A(\myidu/_0079_ ), .Z(\myidu/_0978_ ) );
BUF_X1 \myidu/_1955_ ( .A(\ID_EX_pc [31] ), .Z(\myidu/_0764_ ) );
BUF_X1 \myidu/_1956_ ( .A(\IF_ID_pc [31] ), .Z(\myidu/_0732_ ) );
BUF_X1 \myidu/_1957_ ( .A(\myidu/_0080_ ), .Z(\myidu/_0979_ ) );
BUF_X1 \myidu/_1958_ ( .A(\ID_EX_rs1 [0] ), .Z(\myidu/_0779_ ) );
BUF_X1 \myidu/_1959_ ( .A(\ID_EX_rs1 [1] ), .Z(\myidu/_0780_ ) );
BUF_X1 \myidu/_1960_ ( .A(\ID_EX_rs1 [2] ), .Z(\myidu/_0781_ ) );
BUF_X1 \myidu/_1961_ ( .A(\ID_EX_rs1 [3] ), .Z(\myidu/_0782_ ) );
BUF_X1 \myidu/_1962_ ( .A(\ID_EX_rs1 [4] ), .Z(\myidu/_0783_ ) );
BUF_X1 \myidu/_1963_ ( .A(\ID_EX_rs2 [0] ), .Z(\myidu/_0784_ ) );
BUF_X1 \myidu/_1964_ ( .A(\ID_EX_rs2 [1] ), .Z(\myidu/_0785_ ) );
BUF_X1 \myidu/_1965_ ( .A(\ID_EX_rs2 [2] ), .Z(\myidu/_0786_ ) );
BUF_X1 \myidu/_1966_ ( .A(\ID_EX_rs2 [3] ), .Z(\myidu/_0787_ ) );
BUF_X1 \myidu/_1967_ ( .A(\ID_EX_rs2 [4] ), .Z(\myidu/_0788_ ) );
BUF_X1 \myidu/_1968_ ( .A(\ID_EX_csr [0] ), .Z(\myidu/_0110_ ) );
BUF_X1 \myidu/_1969_ ( .A(\ID_EX_csr [1] ), .Z(\myidu/_0113_ ) );
BUF_X1 \myidu/_1970_ ( .A(\ID_EX_csr [2] ), .Z(\myidu/_0114_ ) );
BUF_X1 \myidu/_1971_ ( .A(\ID_EX_csr [3] ), .Z(\myidu/_0115_ ) );
BUF_X1 \myidu/_1972_ ( .A(\ID_EX_csr [4] ), .Z(\myidu/_0116_ ) );
BUF_X1 \myidu/_1973_ ( .A(\ID_EX_csr [5] ), .Z(\myidu/_0117_ ) );
BUF_X1 \myidu/_1974_ ( .A(\ID_EX_csr [6] ), .Z(\myidu/_0118_ ) );
BUF_X1 \myidu/_1975_ ( .A(\ID_EX_csr [7] ), .Z(\myidu/_0119_ ) );
BUF_X1 \myidu/_1976_ ( .A(\ID_EX_csr [8] ), .Z(\myidu/_0120_ ) );
BUF_X1 \myidu/_1977_ ( .A(\ID_EX_csr [9] ), .Z(\myidu/_0121_ ) );
BUF_X1 \myidu/_1978_ ( .A(\ID_EX_csr [10] ), .Z(\myidu/_0111_ ) );
BUF_X1 \myidu/_1979_ ( .A(\ID_EX_csr [11] ), .Z(\myidu/_0112_ ) );
BUF_X1 \myidu/_1980_ ( .A(stall_quest_loaduse ), .Z(\myidu/_0791_ ) );
BUF_X1 \myidu/_1981_ ( .A(fc_disenable ), .Z(\myidu/_0122_ ) );
BUF_X1 \myidu/_1982_ ( .A(\myidu/_0040_ ), .Z(\myidu/_0939_ ) );
BUF_X1 \myidu/_1983_ ( .A(\myidu/_0041_ ), .Z(\myidu/_0940_ ) );
BUF_X1 \myidu/_1984_ ( .A(\myidu/_0042_ ), .Z(\myidu/_0941_ ) );
BUF_X1 \myidu/_1985_ ( .A(\myidu/_0043_ ), .Z(\myidu/_0942_ ) );
BUF_X1 \myidu/_1986_ ( .A(\myidu/_0044_ ), .Z(\myidu/_0943_ ) );
BUF_X1 \myidu/_1987_ ( .A(\myidu/_0045_ ), .Z(\myidu/_0944_ ) );
BUF_X1 \myidu/_1988_ ( .A(\myidu/_0046_ ), .Z(\myidu/_0945_ ) );
BUF_X1 \myidu/_1989_ ( .A(\myidu/_0047_ ), .Z(\myidu/_0946_ ) );
BUF_X1 \myidu/_1990_ ( .A(\myidu/_0048_ ), .Z(\myidu/_0947_ ) );
BUF_X1 \myidu/_1991_ ( .A(\myidu/_0081_ ), .Z(\myidu/_0980_ ) );
BUF_X1 \myidu/_1992_ ( .A(\myidu/_0082_ ), .Z(\myidu/_0981_ ) );
BUF_X1 \myidu/_1993_ ( .A(\myidu/_0083_ ), .Z(\myidu/_0982_ ) );
BUF_X1 \myidu/_1994_ ( .A(\myidu/_0084_ ), .Z(\myidu/_0983_ ) );
BUF_X1 \myidu/_1995_ ( .A(\myidu/_0085_ ), .Z(\myidu/_0984_ ) );
BUF_X1 \myidu/_1996_ ( .A(\myidu/_0086_ ), .Z(\myidu/_0985_ ) );
BUF_X1 \myidu/_1997_ ( .A(\myidu/_0087_ ), .Z(\myidu/_0986_ ) );
BUF_X1 \myidu/_1998_ ( .A(\myidu/_0088_ ), .Z(\myidu/_0987_ ) );
BUF_X1 \myidu/_1999_ ( .A(\myidu/_0089_ ), .Z(\myidu/_0988_ ) );
BUF_X1 \myidu/_2000_ ( .A(\myidu/_0090_ ), .Z(\myidu/_0989_ ) );
BUF_X1 \myidu/_2001_ ( .A(\myidu/_0091_ ), .Z(\myidu/_0990_ ) );
BUF_X1 \myidu/_2002_ ( .A(\myidu/_0092_ ), .Z(\myidu/_0991_ ) );
BUF_X1 \myidu/_2003_ ( .A(\myidu/_0093_ ), .Z(\myidu/_0992_ ) );
BUF_X1 \myidu/_2004_ ( .A(\myidu/_0094_ ), .Z(\myidu/_0993_ ) );
BUF_X1 \myidu/_2005_ ( .A(\myidu/_0095_ ), .Z(\myidu/_0994_ ) );
BUF_X1 \myidu/_2006_ ( .A(\myidu/_0096_ ), .Z(\myidu/_0995_ ) );
BUF_X1 \myidu/_2007_ ( .A(\myidu/_0097_ ), .Z(\myidu/_0996_ ) );
BUF_X1 \myidu/_2008_ ( .A(\myidu/_0098_ ), .Z(\myidu/_0997_ ) );
BUF_X1 \myidu/_2009_ ( .A(\myidu/_0099_ ), .Z(\myidu/_0998_ ) );
BUF_X1 \myidu/_2010_ ( .A(\myidu/_0100_ ), .Z(\myidu/_0999_ ) );
BUF_X1 \myidu/_2011_ ( .A(\myidu/_0101_ ), .Z(\myidu/_1000_ ) );
BUF_X1 \myidu/_2012_ ( .A(\myidu/_0102_ ), .Z(\myidu/_1001_ ) );
BUF_X1 \myidu/_2013_ ( .A(\myidu/_0103_ ), .Z(\myidu/_1002_ ) );
BUF_X1 \myidu/_2014_ ( .A(\myidu/_0104_ ), .Z(\myidu/_1003_ ) );
BUF_X1 \myidu/_2015_ ( .A(\myidu/_0105_ ), .Z(\myidu/_1004_ ) );
BUF_X1 \myidu/_2016_ ( .A(\myidu/_0106_ ), .Z(\myidu/_1005_ ) );
BUF_X1 \myidu/_2017_ ( .A(\myidu/_0107_ ), .Z(\myidu/_1006_ ) );
BUF_X1 \myidu/_2018_ ( .A(\myidu/_0108_ ), .Z(\myidu/_1007_ ) );
BUF_X1 \myidu/_2019_ ( .A(\myidu/_0109_ ), .Z(\myidu/_1008_ ) );
NOR2_X1 \myifu/_1098_ ( .A1(fanout_net_18 ), .A2(\myifu/_0941_ ), .ZN(\myifu/_0234_ ) );
AND2_X1 \myifu/_1099_ ( .A1(\myifu/_0234_ ), .A2(\myifu/_0942_ ), .ZN(\myifu/_0072_ ) );
INV_X1 \myifu/_1100_ ( .A(\myifu/_0943_ ), .ZN(\myifu/_0235_ ) );
BUF_X4 \myifu/_1101_ ( .A(\myifu/_0235_ ), .Z(\myifu/_0236_ ) );
XNOR2_X1 \myifu/_1102_ ( .A(\myifu/_0888_ ), .B(\myifu/_0063_ ), .ZN(\myifu/_0237_ ) );
XNOR2_X1 \myifu/_1103_ ( .A(\myifu/_0887_ ), .B(\myifu/_0062_ ), .ZN(\myifu/_0238_ ) );
XNOR2_X1 \myifu/_1104_ ( .A(\myifu/_0884_ ), .B(\myifu/_0060_ ), .ZN(\myifu/_0239_ ) );
XNOR2_X1 \myifu/_1105_ ( .A(\myifu/_0885_ ), .B(\myifu/_0061_ ), .ZN(\myifu/_0240_ ) );
AND4_X1 \myifu/_1106_ ( .A1(\myifu/_0237_ ), .A2(\myifu/_0238_ ), .A3(\myifu/_0239_ ), .A4(\myifu/_0240_ ), .ZN(\myifu/_0241_ ) );
XNOR2_X1 \myifu/_1107_ ( .A(\myifu/_0880_ ), .B(\myifu/_0056_ ), .ZN(\myifu/_0242_ ) );
XNOR2_X1 \myifu/_1108_ ( .A(\myifu/_0881_ ), .B(\myifu/_0057_ ), .ZN(\myifu/_0243_ ) );
XNOR2_X1 \myifu/_1109_ ( .A(\myifu/_0882_ ), .B(\myifu/_0058_ ), .ZN(\myifu/_0244_ ) );
XNOR2_X1 \myifu/_1110_ ( .A(\myifu/_0883_ ), .B(\myifu/_0059_ ), .ZN(\myifu/_0245_ ) );
AND4_X1 \myifu/_1111_ ( .A1(\myifu/_0242_ ), .A2(\myifu/_0243_ ), .A3(\myifu/_0244_ ), .A4(\myifu/_0245_ ), .ZN(\myifu/_0246_ ) );
XNOR2_X1 \myifu/_1112_ ( .A(\myifu/_0877_ ), .B(\myifu/_0053_ ), .ZN(\myifu/_0247_ ) );
XNOR2_X1 \myifu/_1113_ ( .A(\myifu/_0878_ ), .B(\myifu/_0054_ ), .ZN(\myifu/_0248_ ) );
XNOR2_X1 \myifu/_1114_ ( .A(\myifu/_0879_ ), .B(\myifu/_0055_ ), .ZN(\myifu/_0249_ ) );
XNOR2_X1 \myifu/_1115_ ( .A(\myifu/_0876_ ), .B(\myifu/_0052_ ), .ZN(\myifu/_0250_ ) );
AND4_X1 \myifu/_1116_ ( .A1(\myifu/_0247_ ), .A2(\myifu/_0248_ ), .A3(\myifu/_0249_ ), .A4(\myifu/_0250_ ), .ZN(\myifu/_0251_ ) );
XNOR2_X1 \myifu/_1117_ ( .A(\myifu/_0872_ ), .B(\myifu/_0049_ ), .ZN(\myifu/_0252_ ) );
XNOR2_X1 \myifu/_1118_ ( .A(\myifu/_0874_ ), .B(\myifu/_0051_ ), .ZN(\myifu/_0253_ ) );
XNOR2_X1 \myifu/_1119_ ( .A(\myifu/_0873_ ), .B(\myifu/_0050_ ), .ZN(\myifu/_0254_ ) );
XNOR2_X1 \myifu/_1120_ ( .A(\myifu/_0871_ ), .B(\myifu/_0048_ ), .ZN(\myifu/_0255_ ) );
AND4_X1 \myifu/_1121_ ( .A1(\myifu/_0252_ ), .A2(\myifu/_0253_ ), .A3(\myifu/_0254_ ), .A4(\myifu/_0255_ ), .ZN(\myifu/_0256_ ) );
AND4_X1 \myifu/_1122_ ( .A1(\myifu/_0241_ ), .A2(\myifu/_0246_ ), .A3(\myifu/_0251_ ), .A4(\myifu/_0256_ ), .ZN(\myifu/_0257_ ) );
XNOR2_X1 \myifu/_1123_ ( .A(\myifu/_0864_ ), .B(\myifu/_0861_ ), .ZN(\myifu/_0258_ ) );
XNOR2_X1 \myifu/_1124_ ( .A(\myifu/_0893_ ), .B(\myifu/_0068_ ), .ZN(\myifu/_0259_ ) );
XNOR2_X1 \myifu/_1125_ ( .A(\myifu/_0892_ ), .B(\myifu/_0067_ ), .ZN(\myifu/_0260_ ) );
XNOR2_X1 \myifu/_1126_ ( .A(\myifu/_0890_ ), .B(\myifu/_0065_ ), .ZN(\myifu/_0261_ ) );
XNOR2_X1 \myifu/_1127_ ( .A(\myifu/_0891_ ), .B(\myifu/_0066_ ), .ZN(\myifu/_0262_ ) );
AND4_X1 \myifu/_1128_ ( .A1(\myifu/_0259_ ), .A2(\myifu/_0260_ ), .A3(\myifu/_0261_ ), .A4(\myifu/_0262_ ), .ZN(\myifu/_0263_ ) );
XNOR2_X1 \myifu/_1129_ ( .A(\myifu/_0875_ ), .B(\myifu/_0862_ ), .ZN(\myifu/_0264_ ) );
XOR2_X1 \myifu/_1130_ ( .A(\myifu/_0886_ ), .B(\myifu/_0863_ ), .Z(\myifu/_0265_ ) );
INV_X1 \myifu/_1131_ ( .A(\myifu/_0064_ ), .ZN(\myifu/_0266_ ) );
AND2_X1 \myifu/_1132_ ( .A1(\myifu/_0266_ ), .A2(\myifu/_0889_ ), .ZN(\myifu/_0267_ ) );
NOR2_X1 \myifu/_1133_ ( .A1(\myifu/_0266_ ), .A2(\myifu/_0889_ ), .ZN(\myifu/_0268_ ) );
NOR3_X1 \myifu/_1134_ ( .A1(\myifu/_0265_ ), .A2(\myifu/_0267_ ), .A3(\myifu/_0268_ ), .ZN(\myifu/_0269_ ) );
AND4_X1 \myifu/_1135_ ( .A1(\myifu/_0258_ ), .A2(\myifu/_0263_ ), .A3(\myifu/_0264_ ), .A4(\myifu/_0269_ ), .ZN(\myifu/_0270_ ) );
XNOR2_X1 \myifu/_1136_ ( .A(\myifu/_0867_ ), .B(\myifu/_0044_ ), .ZN(\myifu/_0271_ ) );
XNOR2_X1 \myifu/_1137_ ( .A(\myifu/_0870_ ), .B(\myifu/_0047_ ), .ZN(\myifu/_0272_ ) );
XNOR2_X1 \myifu/_1138_ ( .A(\myifu/_0869_ ), .B(\myifu/_0046_ ), .ZN(\myifu/_0273_ ) );
XNOR2_X1 \myifu/_1139_ ( .A(\myifu/_0868_ ), .B(\myifu/_0045_ ), .ZN(\myifu/_0274_ ) );
AND4_X1 \myifu/_1140_ ( .A1(\myifu/_0271_ ), .A2(\myifu/_0272_ ), .A3(\myifu/_0273_ ), .A4(\myifu/_0274_ ), .ZN(\myifu/_0275_ ) );
XNOR2_X1 \myifu/_1141_ ( .A(\myifu/_0894_ ), .B(\myifu/_0069_ ), .ZN(\myifu/_0276_ ) );
XNOR2_X1 \myifu/_1142_ ( .A(\myifu/_0895_ ), .B(\myifu/_0070_ ), .ZN(\myifu/_0277_ ) );
XNOR2_X1 \myifu/_1143_ ( .A(\myifu/_0865_ ), .B(\myifu/_0042_ ), .ZN(\myifu/_0278_ ) );
XNOR2_X1 \myifu/_1144_ ( .A(\myifu/_0866_ ), .B(\myifu/_0043_ ), .ZN(\myifu/_0279_ ) );
AND4_X1 \myifu/_1145_ ( .A1(\myifu/_0276_ ), .A2(\myifu/_0277_ ), .A3(\myifu/_0278_ ), .A4(\myifu/_0279_ ), .ZN(\myifu/_0280_ ) );
NAND4_X1 \myifu/_1146_ ( .A1(\myifu/_0257_ ), .A2(\myifu/_0270_ ), .A3(\myifu/_0275_ ), .A4(\myifu/_0280_ ), .ZN(\myifu/_0281_ ) );
AOI21_X1 \myifu/_1147_ ( .A(\myifu/_0236_ ), .B1(\myifu/_0281_ ), .B2(\myifu/_0141_ ), .ZN(\myifu/_0973_ ) );
INV_X1 \myifu/_1148_ ( .A(\myifu/_0234_ ), .ZN(\myifu/_0025_ ) );
INV_X1 \myifu/_1149_ ( .A(\myifu/_0067_ ), .ZN(\myifu/_0282_ ) );
NOR2_X1 \myifu/_1150_ ( .A1(\myifu/_0282_ ), .A2(\myifu/_0956_ ), .ZN(\myifu/_0283_ ) );
INV_X1 \myifu/_1151_ ( .A(\myifu/_0046_ ), .ZN(\myifu/_0284_ ) );
INV_X1 \myifu/_1152_ ( .A(\myifu/_0058_ ), .ZN(\myifu/_0285_ ) );
OAI22_X1 \myifu/_1153_ ( .A1(\myifu/_0284_ ), .A2(\myifu/_0971_ ), .B1(\myifu/_0285_ ), .B2(\myifu/_0958_ ), .ZN(\myifu/_0286_ ) );
AOI211_X4 \myifu/_1154_ ( .A(\myifu/_0283_ ), .B(\myifu/_0286_ ), .C1(\myifu/_0284_ ), .C2(\myifu/_0971_ ), .ZN(\myifu/_0287_ ) );
INV_X1 \myifu/_1155_ ( .A(\myifu/_0055_ ), .ZN(\myifu/_0288_ ) );
AOI22_X1 \myifu/_1156_ ( .A1(\myifu/_0288_ ), .A2(\myifu/_0954_ ), .B1(\myifu/_0285_ ), .B2(\myifu/_0958_ ), .ZN(\myifu/_0289_ ) );
AND2_X1 \myifu/_1157_ ( .A1(\myifu/_0053_ ), .A2(\myifu/_0952_ ), .ZN(\myifu/_0290_ ) );
NOR2_X1 \myifu/_1158_ ( .A1(\myifu/_0053_ ), .A2(\myifu/_0952_ ), .ZN(\myifu/_0291_ ) );
OAI211_X2 \myifu/_1159_ ( .A(\myifu/_0287_ ), .B(\myifu/_0289_ ), .C1(\myifu/_0290_ ), .C2(\myifu/_0291_ ), .ZN(\myifu/_0292_ ) );
INV_X1 \myifu/_1160_ ( .A(\myifu/_0066_ ), .ZN(\myifu/_0293_ ) );
INV_X1 \myifu/_1161_ ( .A(\myifu/_0048_ ), .ZN(\myifu/_0294_ ) );
AOI22_X1 \myifu/_1162_ ( .A1(\myifu/_0293_ ), .A2(\myifu/_0945_ ), .B1(\myifu/_0294_ ), .B2(\myifu/_0947_ ), .ZN(\myifu/_0295_ ) );
INV_X1 \myifu/_1163_ ( .A(\myifu/_0966_ ), .ZN(\myifu/_0296_ ) );
OAI221_X1 \myifu/_1164_ ( .A(\myifu/_0295_ ), .B1(\myifu/_0293_ ), .B2(\myifu/_0945_ ), .C1(\myifu/_0070_ ), .C2(\myifu/_0296_ ), .ZN(\myifu/_0297_ ) );
INV_X1 \myifu/_1165_ ( .A(\myifu/_0043_ ), .ZN(\myifu/_0298_ ) );
AOI22_X1 \myifu/_1166_ ( .A1(\myifu/_0070_ ), .A2(\myifu/_0296_ ), .B1(\myifu/_0298_ ), .B2(\myifu/_0968_ ), .ZN(\myifu/_0299_ ) );
INV_X1 \myifu/_1167_ ( .A(\myifu/_0047_ ), .ZN(\myifu/_0300_ ) );
NAND2_X1 \myifu/_1168_ ( .A1(\myifu/_0300_ ), .A2(\myifu/_0946_ ), .ZN(\myifu/_0301_ ) );
OAI211_X2 \myifu/_1169_ ( .A(\myifu/_0299_ ), .B(\myifu/_0301_ ), .C1(\myifu/_0298_ ), .C2(\myifu/_0968_ ), .ZN(\myifu/_0302_ ) );
NOR3_X1 \myifu/_1170_ ( .A1(\myifu/_0292_ ), .A2(\myifu/_0297_ ), .A3(\myifu/_0302_ ), .ZN(\myifu/_0303_ ) );
XNOR2_X1 \myifu/_1171_ ( .A(\myifu/_0045_ ), .B(\myifu/_0970_ ), .ZN(\myifu/_0304_ ) );
INV_X1 \myifu/_1172_ ( .A(\myifu/_0069_ ), .ZN(\myifu/_0305_ ) );
INV_X1 \myifu/_1173_ ( .A(\myifu/_0052_ ), .ZN(\myifu/_0306_ ) );
OAI221_X1 \myifu/_1174_ ( .A(\myifu/_0304_ ), .B1(\myifu/_0305_ ), .B2(\myifu/_0965_ ), .C1(\myifu/_0306_ ), .C2(\myifu/_0951_ ), .ZN(\myifu/_0307_ ) );
XOR2_X1 \myifu/_1175_ ( .A(\myifu/_0049_ ), .B(\myifu/_0948_ ), .Z(\myifu/_0308_ ) );
XOR2_X1 \myifu/_1176_ ( .A(\myifu/_0068_ ), .B(\myifu/_0964_ ), .Z(\myifu/_0309_ ) );
NOR3_X1 \myifu/_1177_ ( .A1(\myifu/_0307_ ), .A2(\myifu/_0308_ ), .A3(\myifu/_0309_ ), .ZN(\myifu/_0310_ ) );
INV_X1 \myifu/_1178_ ( .A(\myifu/_0044_ ), .ZN(\myifu/_0311_ ) );
INV_X1 \myifu/_1179_ ( .A(\myifu/_0054_ ), .ZN(\myifu/_0312_ ) );
OAI22_X1 \myifu/_1180_ ( .A1(\myifu/_0311_ ), .A2(\myifu/_0969_ ), .B1(\myifu/_0312_ ), .B2(\myifu/_0953_ ), .ZN(\myifu/_0313_ ) );
XNOR2_X1 \myifu/_1181_ ( .A(\myifu/_0051_ ), .B(\myifu/_0950_ ), .ZN(\myifu/_0314_ ) );
INV_X1 \myifu/_1182_ ( .A(\myifu/_0050_ ), .ZN(\myifu/_0315_ ) );
OAI221_X1 \myifu/_1183_ ( .A(\myifu/_0314_ ), .B1(\myifu/_0315_ ), .B2(\myifu/_0949_ ), .C1(\myifu/_0288_ ), .C2(\myifu/_0954_ ), .ZN(\myifu/_0316_ ) );
AOI211_X4 \myifu/_1184_ ( .A(\myifu/_0313_ ), .B(\myifu/_0316_ ), .C1(\myifu/_0315_ ), .C2(\myifu/_0949_ ), .ZN(\myifu/_0317_ ) );
AND3_X1 \myifu/_1185_ ( .A1(\myifu/_0303_ ), .A2(\myifu/_0310_ ), .A3(\myifu/_0317_ ), .ZN(\myifu/_0318_ ) );
OAI22_X1 \myifu/_1186_ ( .A1(\myifu/_0300_ ), .A2(\myifu/_0946_ ), .B1(\myifu/_0294_ ), .B2(\myifu/_0947_ ), .ZN(\myifu/_0319_ ) );
AOI221_X4 \myifu/_1187_ ( .A(\myifu/_0319_ ), .B1(\myifu/_0305_ ), .B2(\myifu/_0965_ ), .C1(\myifu/_0311_ ), .C2(\myifu/_0969_ ), .ZN(\myifu/_0320_ ) );
XNOR2_X1 \myifu/_1188_ ( .A(\myifu/_0057_ ), .B(\myifu/_0957_ ), .ZN(\myifu/_0321_ ) );
INV_X1 \myifu/_1189_ ( .A(\myifu/_0063_ ), .ZN(\myifu/_0322_ ) );
NAND2_X1 \myifu/_1190_ ( .A1(\myifu/_0322_ ), .A2(\myifu/_0963_ ), .ZN(\myifu/_0323_ ) );
NAND4_X1 \myifu/_1191_ ( .A1(\myifu/_0320_ ), .A2(\myifu/_0975_ ), .A3(\myifu/_0321_ ), .A4(\myifu/_0323_ ), .ZN(\myifu/_0324_ ) );
INV_X1 \myifu/_1192_ ( .A(\myifu/_0955_ ), .ZN(\myifu/_0325_ ) );
AOI22_X1 \myifu/_1193_ ( .A1(\myifu/_0282_ ), .A2(\myifu/_0956_ ), .B1(\myifu/_0325_ ), .B2(\myifu/_0056_ ), .ZN(\myifu/_0326_ ) );
NAND2_X1 \myifu/_1194_ ( .A1(\myifu/_0306_ ), .A2(\myifu/_0951_ ), .ZN(\myifu/_0327_ ) );
INV_X1 \myifu/_1195_ ( .A(\myifu/_0061_ ), .ZN(\myifu/_0328_ ) );
OAI211_X2 \myifu/_1196_ ( .A(\myifu/_0326_ ), .B(\myifu/_0327_ ), .C1(\myifu/_0328_ ), .C2(\myifu/_0961_ ), .ZN(\myifu/_0329_ ) );
XOR2_X1 \myifu/_1197_ ( .A(\myifu/_0059_ ), .B(\myifu/_0959_ ), .Z(\myifu/_0330_ ) );
OAI22_X1 \myifu/_1198_ ( .A1(\myifu/_0056_ ), .A2(\myifu/_0325_ ), .B1(\myifu/_0322_ ), .B2(\myifu/_0963_ ), .ZN(\myifu/_0331_ ) );
OR3_X1 \myifu/_1199_ ( .A1(\myifu/_0329_ ), .A2(\myifu/_0330_ ), .A3(\myifu/_0331_ ), .ZN(\myifu/_0332_ ) );
INV_X1 \myifu/_1200_ ( .A(\myifu/_0060_ ), .ZN(\myifu/_0333_ ) );
INV_X1 \myifu/_1201_ ( .A(\myifu/_0062_ ), .ZN(\myifu/_0334_ ) );
AOI22_X1 \myifu/_1202_ ( .A1(\myifu/_0333_ ), .A2(\myifu/_0960_ ), .B1(\myifu/_0334_ ), .B2(\myifu/_0962_ ), .ZN(\myifu/_0335_ ) );
NAND2_X1 \myifu/_1203_ ( .A1(\myifu/_0328_ ), .A2(\myifu/_0961_ ), .ZN(\myifu/_0336_ ) );
OAI211_X2 \myifu/_1204_ ( .A(\myifu/_0335_ ), .B(\myifu/_0336_ ), .C1(\myifu/_0334_ ), .C2(\myifu/_0962_ ), .ZN(\myifu/_0337_ ) );
INV_X1 \myifu/_1205_ ( .A(\myifu/_0042_ ), .ZN(\myifu/_0338_ ) );
AOI22_X1 \myifu/_1206_ ( .A1(\myifu/_0338_ ), .A2(\myifu/_0967_ ), .B1(\myifu/_0312_ ), .B2(\myifu/_0953_ ), .ZN(\myifu/_0339_ ) );
OAI221_X1 \myifu/_1207_ ( .A(\myifu/_0339_ ), .B1(\myifu/_0338_ ), .B2(\myifu/_0967_ ), .C1(\myifu/_0333_ ), .C2(\myifu/_0960_ ), .ZN(\myifu/_0340_ ) );
NOR4_X1 \myifu/_1208_ ( .A1(\myifu/_0324_ ), .A2(\myifu/_0332_ ), .A3(\myifu/_0337_ ), .A4(\myifu/_0340_ ), .ZN(\myifu/_0341_ ) );
NAND3_X1 \myifu/_1209_ ( .A1(\myifu/_0318_ ), .A2(\myifu/_0072_ ), .A3(\myifu/_0341_ ), .ZN(\myifu/_0342_ ) );
INV_X1 \myifu/_1210_ ( .A(fanout_net_18 ), .ZN(\myifu/_0343_ ) );
INV_X1 \myifu/_1211_ ( .A(\myifu/_0929_ ), .ZN(\myifu/_0344_ ) );
BUF_X4 \myifu/_1212_ ( .A(\myifu/_0344_ ), .Z(\myifu/_0345_ ) );
NAND3_X1 \myifu/_1213_ ( .A1(\myifu/_0343_ ), .A2(\myifu/_0345_ ), .A3(\myifu/_0943_ ), .ZN(\myifu/_0346_ ) );
OR3_X1 \myifu/_1214_ ( .A1(\myifu/_0938_ ), .A2(\myifu/_0932_ ), .A3(\myifu/_0934_ ), .ZN(\myifu/_0347_ ) );
INV_X1 \myifu/_1215_ ( .A(\myifu/_0939_ ), .ZN(\myifu/_0348_ ) );
INV_X1 \myifu/_1216_ ( .A(\myifu/_0933_ ), .ZN(\myifu/_0349_ ) );
NAND4_X1 \myifu/_1217_ ( .A1(\myifu/_0348_ ), .A2(\myifu/_0349_ ), .A3(\myifu/_0940_ ), .A4(\myifu/_0931_ ), .ZN(\myifu/_0350_ ) );
NOR2_X1 \myifu/_1218_ ( .A1(\myifu/_0347_ ), .A2(\myifu/_0350_ ), .ZN(\myifu/_0351_ ) );
CLKBUF_X2 \myifu/_1219_ ( .A(\myifu/_0351_ ), .Z(\myifu/_0352_ ) );
NAND4_X1 \myifu/_1220_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0343_ ), .A3(\myifu/_0935_ ), .A4(fanout_net_19 ), .ZN(\myifu/_0353_ ) );
NAND3_X1 \myifu/_1221_ ( .A1(\myifu/_0342_ ), .A2(\myifu/_0346_ ), .A3(\myifu/_0353_ ), .ZN(\myifu/_0022_ ) );
AND2_X1 \myifu/_1222_ ( .A1(\myifu/_0318_ ), .A2(\myifu/_0341_ ), .ZN(\myifu/_0354_ ) );
INV_X1 \myifu/_1223_ ( .A(\myifu/_0354_ ), .ZN(\myifu/_0355_ ) );
NAND3_X1 \myifu/_1224_ ( .A1(\myifu/_0355_ ), .A2(\myifu/_0071_ ), .A3(\myifu/_0072_ ), .ZN(\myifu/_0356_ ) );
AND2_X1 \myifu/_1225_ ( .A1(\myifu/_0351_ ), .A2(\myifu/_0935_ ), .ZN(\myifu/_0357_ ) );
INV_X2 \myifu/_1226_ ( .A(fanout_net_19 ), .ZN(\myifu/_0358_ ) );
OR3_X1 \myifu/_1227_ ( .A1(\myifu/_0357_ ), .A2(fanout_net_18 ), .A3(\myifu/_0358_ ), .ZN(\myifu/_0359_ ) );
NAND2_X1 \myifu/_1228_ ( .A1(\myifu/_0356_ ), .A2(\myifu/_0359_ ), .ZN(\myifu/_0023_ ) );
INV_X1 \myifu/_1229_ ( .A(\myifu/_0072_ ), .ZN(\myifu/_0360_ ) );
NOR3_X1 \myifu/_1230_ ( .A1(\myifu/_0354_ ), .A2(\myifu/_0071_ ), .A3(\myifu/_0360_ ), .ZN(\myifu/_0361_ ) );
AND2_X1 \myifu/_1231_ ( .A1(\myifu/_0943_ ), .A2(\myifu/_0929_ ), .ZN(\myifu/_0362_ ) );
AND2_X1 \myifu/_1232_ ( .A1(\myifu/_0941_ ), .A2(\myifu/_0942_ ), .ZN(\myifu/_0363_ ) );
OR4_X1 \myifu/_1233_ ( .A1(fanout_net_18 ), .A2(\myifu/_0361_ ), .A3(\myifu/_0362_ ), .A4(\myifu/_0363_ ), .ZN(\myifu/_0021_ ) );
BUF_X4 \myifu/_1234_ ( .A(\myifu/_0358_ ), .Z(\myifu/_0364_ ) );
OAI21_X1 \myifu/_1235_ ( .A(\myifu/_0364_ ), .B1(\myifu/_0354_ ), .B2(\myifu/_0360_ ), .ZN(\myifu/_0937_ ) );
INV_X1 \myifu/_1236_ ( .A(\myifu/_0942_ ), .ZN(\myifu/_0365_ ) );
OAI21_X1 \myifu/_1237_ ( .A(\myifu/_0364_ ), .B1(\myifu/_0354_ ), .B2(\myifu/_0365_ ), .ZN(\myifu/_0936_ ) );
INV_X1 \myifu/_1238_ ( .A(\myifu/_0861_ ), .ZN(\myifu/_0366_ ) );
NOR2_X1 \myifu/_1239_ ( .A1(\myifu/_0366_ ), .A2(\myifu/_0974_ ), .ZN(\myifu/_0858_ ) );
INV_X1 \myifu/_1240_ ( .A(\myifu/_0862_ ), .ZN(\myifu/_0367_ ) );
NOR2_X1 \myifu/_1241_ ( .A1(\myifu/_0367_ ), .A2(\myifu/_0974_ ), .ZN(\myifu/_0859_ ) );
MUX2_X1 \myifu/_1242_ ( .A(\myifu/_0863_ ), .B(\myifu/_0972_ ), .S(\myifu/_0974_ ), .Z(\myifu/_0860_ ) );
NOR2_X1 \myifu/_1243_ ( .A1(\myifu/_0942_ ), .A2(fanout_net_19 ), .ZN(\myifu/_0368_ ) );
NOR2_X1 \myifu/_1244_ ( .A1(\myifu/_0363_ ), .A2(\myifu/_0368_ ), .ZN(\myifu/_0369_ ) );
OAI21_X1 \myifu/_1245_ ( .A(\myifu/_0369_ ), .B1(\myifu/_0354_ ), .B2(\myifu/_0365_ ), .ZN(\myifu/_0370_ ) );
OR2_X2 \myifu/_1246_ ( .A1(\myifu/_0370_ ), .A2(fanout_net_18 ), .ZN(\myifu/_0371_ ) );
BUF_X4 \myifu/_1247_ ( .A(\myifu/_0371_ ), .Z(\myifu/_0372_ ) );
INV_X1 \myifu/_1248_ ( .A(\myifu/_0972_ ), .ZN(\myifu/_0373_ ) );
OAI211_X2 \myifu/_1249_ ( .A(\myifu/_0367_ ), .B(\myifu/_0026_ ), .C1(\myifu/_0373_ ), .C2(\myifu/_0863_ ), .ZN(\myifu/_0374_ ) );
INV_X1 \myifu/_1250_ ( .A(\myifu/_0863_ ), .ZN(\myifu/_0375_ ) );
NOR2_X1 \myifu/_1251_ ( .A1(\myifu/_0375_ ), .A2(\myifu/_0972_ ), .ZN(\myifu/_0376_ ) );
NOR2_X1 \myifu/_1252_ ( .A1(\myifu/_0374_ ), .A2(\myifu/_0376_ ), .ZN(\myifu/_0377_ ) );
AOI21_X2 \myifu/_1253_ ( .A(\myifu/_0358_ ), .B1(\myifu/_0351_ ), .B2(\myifu/_0377_ ), .ZN(\myifu/_0378_ ) );
BUF_X4 \myifu/_1254_ ( .A(\myifu/_0378_ ), .Z(\myifu/_0379_ ) );
OAI21_X1 \myifu/_1255_ ( .A(\myifu/_0174_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0380_ ) );
NOR2_X2 \myifu/_1256_ ( .A1(\myifu/_0370_ ), .A2(fanout_net_18 ), .ZN(\myifu/_0381_ ) );
BUF_X8 \myifu/_1257_ ( .A(\myifu/_0381_ ), .Z(\myifu/_0382_ ) );
OR2_X1 \myifu/_1258_ ( .A1(fanout_net_19 ), .A2(\myifu/_0142_ ), .ZN(\myifu/_0383_ ) );
CLKBUF_X2 \myifu/_1259_ ( .A(\myifu/_0377_ ), .Z(\myifu/_0384_ ) );
AND3_X1 \myifu/_1260_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0897_ ), .ZN(\myifu/_0385_ ) );
OAI211_X2 \myifu/_1261_ ( .A(\myifu/_0382_ ), .B(\myifu/_0383_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0385_ ), .ZN(\myifu/_0386_ ) );
NAND2_X1 \myifu/_1262_ ( .A1(\myifu/_0380_ ), .A2(\myifu/_0386_ ), .ZN(\myifu/_0106_ ) );
OAI21_X1 \myifu/_1263_ ( .A(\myifu/_0185_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0387_ ) );
OR2_X1 \myifu/_1264_ ( .A1(fanout_net_19 ), .A2(\myifu/_0153_ ), .ZN(\myifu/_0388_ ) );
AND3_X1 \myifu/_1265_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0908_ ), .ZN(\myifu/_0389_ ) );
OAI211_X2 \myifu/_1266_ ( .A(\myifu/_0382_ ), .B(\myifu/_0388_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0389_ ), .ZN(\myifu/_0390_ ) );
NAND2_X1 \myifu/_1267_ ( .A1(\myifu/_0387_ ), .A2(\myifu/_0390_ ), .ZN(\myifu/_0107_ ) );
OAI21_X1 \myifu/_1268_ ( .A(\myifu/_0196_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0391_ ) );
OR2_X1 \myifu/_1269_ ( .A1(fanout_net_19 ), .A2(\myifu/_0164_ ), .ZN(\myifu/_0392_ ) );
AND3_X1 \myifu/_1270_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0919_ ), .ZN(\myifu/_0393_ ) );
OAI211_X2 \myifu/_1271_ ( .A(\myifu/_0382_ ), .B(\myifu/_0392_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0393_ ), .ZN(\myifu/_0394_ ) );
NAND2_X1 \myifu/_1272_ ( .A1(\myifu/_0391_ ), .A2(\myifu/_0394_ ), .ZN(\myifu/_0108_ ) );
OAI21_X1 \myifu/_1273_ ( .A(\myifu/_0198_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0395_ ) );
OR2_X1 \myifu/_1274_ ( .A1(fanout_net_19 ), .A2(\myifu/_0167_ ), .ZN(\myifu/_0396_ ) );
AND3_X1 \myifu/_1275_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0922_ ), .ZN(\myifu/_0397_ ) );
OAI211_X2 \myifu/_1276_ ( .A(\myifu/_0382_ ), .B(\myifu/_0396_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0397_ ), .ZN(\myifu/_0398_ ) );
NAND2_X1 \myifu/_1277_ ( .A1(\myifu/_0395_ ), .A2(\myifu/_0398_ ), .ZN(\myifu/_0109_ ) );
OAI21_X1 \myifu/_1278_ ( .A(\myifu/_0199_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0399_ ) );
OR2_X1 \myifu/_1279_ ( .A1(fanout_net_19 ), .A2(\myifu/_0168_ ), .ZN(\myifu/_0400_ ) );
AND3_X1 \myifu/_1280_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0923_ ), .ZN(\myifu/_0401_ ) );
OAI211_X2 \myifu/_1281_ ( .A(\myifu/_0382_ ), .B(\myifu/_0400_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0401_ ), .ZN(\myifu/_0402_ ) );
NAND2_X1 \myifu/_1282_ ( .A1(\myifu/_0399_ ), .A2(\myifu/_0402_ ), .ZN(\myifu/_0110_ ) );
OAI21_X1 \myifu/_1283_ ( .A(\myifu/_0200_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0403_ ) );
OR2_X1 \myifu/_1284_ ( .A1(fanout_net_19 ), .A2(\myifu/_0169_ ), .ZN(\myifu/_0404_ ) );
AND3_X1 \myifu/_1285_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0924_ ), .ZN(\myifu/_0405_ ) );
OAI211_X2 \myifu/_1286_ ( .A(\myifu/_0382_ ), .B(\myifu/_0404_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0405_ ), .ZN(\myifu/_0406_ ) );
NAND2_X1 \myifu/_1287_ ( .A1(\myifu/_0403_ ), .A2(\myifu/_0406_ ), .ZN(\myifu/_0111_ ) );
OAI21_X1 \myifu/_1288_ ( .A(\myifu/_0201_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0407_ ) );
OR2_X1 \myifu/_1289_ ( .A1(fanout_net_19 ), .A2(\myifu/_0170_ ), .ZN(\myifu/_0408_ ) );
AND3_X1 \myifu/_1290_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0925_ ), .ZN(\myifu/_0409_ ) );
OAI211_X2 \myifu/_1291_ ( .A(\myifu/_0382_ ), .B(\myifu/_0408_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0409_ ), .ZN(\myifu/_0410_ ) );
NAND2_X1 \myifu/_1292_ ( .A1(\myifu/_0407_ ), .A2(\myifu/_0410_ ), .ZN(\myifu/_0112_ ) );
OAI21_X1 \myifu/_1293_ ( .A(\myifu/_0202_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0411_ ) );
OR2_X1 \myifu/_1294_ ( .A1(fanout_net_19 ), .A2(\myifu/_0171_ ), .ZN(\myifu/_0412_ ) );
AND3_X1 \myifu/_1295_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0926_ ), .ZN(\myifu/_0413_ ) );
OAI211_X2 \myifu/_1296_ ( .A(\myifu/_0382_ ), .B(\myifu/_0412_ ), .C1(\myifu/_0364_ ), .C2(\myifu/_0413_ ), .ZN(\myifu/_0414_ ) );
NAND2_X1 \myifu/_1297_ ( .A1(\myifu/_0411_ ), .A2(\myifu/_0414_ ), .ZN(\myifu/_0113_ ) );
OAI21_X1 \myifu/_1298_ ( .A(\myifu/_0203_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0415_ ) );
OR2_X1 \myifu/_1299_ ( .A1(fanout_net_19 ), .A2(\myifu/_0172_ ), .ZN(\myifu/_0416_ ) );
BUF_X4 \myifu/_1300_ ( .A(\myifu/_0358_ ), .Z(\myifu/_0417_ ) );
AND3_X1 \myifu/_1301_ ( .A1(\myifu/_0352_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0927_ ), .ZN(\myifu/_0418_ ) );
OAI211_X2 \myifu/_1302_ ( .A(\myifu/_0382_ ), .B(\myifu/_0416_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0418_ ), .ZN(\myifu/_0419_ ) );
NAND2_X1 \myifu/_1303_ ( .A1(\myifu/_0415_ ), .A2(\myifu/_0419_ ), .ZN(\myifu/_0114_ ) );
OAI21_X1 \myifu/_1304_ ( .A(\myifu/_0204_ ), .B1(\myifu/_0372_ ), .B2(\myifu/_0379_ ), .ZN(\myifu/_0420_ ) );
OR2_X1 \myifu/_1305_ ( .A1(fanout_net_19 ), .A2(\myifu/_0173_ ), .ZN(\myifu/_0421_ ) );
CLKBUF_X2 \myifu/_1306_ ( .A(\myifu/_0351_ ), .Z(\myifu/_0422_ ) );
AND3_X1 \myifu/_1307_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0384_ ), .A3(\myifu/_0928_ ), .ZN(\myifu/_0423_ ) );
OAI211_X2 \myifu/_1308_ ( .A(\myifu/_0382_ ), .B(\myifu/_0421_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0423_ ), .ZN(\myifu/_0424_ ) );
NAND2_X1 \myifu/_1309_ ( .A1(\myifu/_0420_ ), .A2(\myifu/_0424_ ), .ZN(\myifu/_0115_ ) );
BUF_X4 \myifu/_1310_ ( .A(\myifu/_0371_ ), .Z(\myifu/_0425_ ) );
BUF_X4 \myifu/_1311_ ( .A(\myifu/_0378_ ), .Z(\myifu/_0426_ ) );
OAI21_X1 \myifu/_1312_ ( .A(\myifu/_0175_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0427_ ) );
BUF_X8 \myifu/_1313_ ( .A(\myifu/_0381_ ), .Z(\myifu/_0428_ ) );
OR2_X1 \myifu/_1314_ ( .A1(fanout_net_19 ), .A2(\myifu/_0143_ ), .ZN(\myifu/_0429_ ) );
CLKBUF_X2 \myifu/_1315_ ( .A(\myifu/_0377_ ), .Z(\myifu/_0430_ ) );
AND3_X1 \myifu/_1316_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0898_ ), .ZN(\myifu/_0431_ ) );
OAI211_X2 \myifu/_1317_ ( .A(\myifu/_0428_ ), .B(\myifu/_0429_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0431_ ), .ZN(\myifu/_0432_ ) );
NAND2_X1 \myifu/_1318_ ( .A1(\myifu/_0427_ ), .A2(\myifu/_0432_ ), .ZN(\myifu/_0116_ ) );
OAI21_X1 \myifu/_1319_ ( .A(\myifu/_0176_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0433_ ) );
OR2_X1 \myifu/_1320_ ( .A1(fanout_net_19 ), .A2(\myifu/_0144_ ), .ZN(\myifu/_0434_ ) );
AND3_X1 \myifu/_1321_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0899_ ), .ZN(\myifu/_0435_ ) );
OAI211_X2 \myifu/_1322_ ( .A(\myifu/_0428_ ), .B(\myifu/_0434_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0435_ ), .ZN(\myifu/_0436_ ) );
NAND2_X1 \myifu/_1323_ ( .A1(\myifu/_0433_ ), .A2(\myifu/_0436_ ), .ZN(\myifu/_0117_ ) );
BUF_X8 \myifu/_1324_ ( .A(\myifu/_0381_ ), .Z(\myifu/_0437_ ) );
OR2_X1 \myifu/_1325_ ( .A1(fanout_net_19 ), .A2(\myifu/_0145_ ), .ZN(\myifu/_0438_ ) );
BUF_X4 \myifu/_1326_ ( .A(\myifu/_0358_ ), .Z(\myifu/_0439_ ) );
CLKBUF_X2 \myifu/_1327_ ( .A(\myifu/_0351_ ), .Z(\myifu/_0440_ ) );
CLKBUF_X2 \myifu/_1328_ ( .A(\myifu/_0377_ ), .Z(\myifu/_0441_ ) );
AND3_X1 \myifu/_1329_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0900_ ), .ZN(\myifu/_0442_ ) );
OAI211_X2 \myifu/_1330_ ( .A(\myifu/_0437_ ), .B(\myifu/_0438_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0442_ ), .ZN(\myifu/_0443_ ) );
NOR2_X1 \myifu/_1331_ ( .A1(\myifu/_0371_ ), .A2(\myifu/_0378_ ), .ZN(\myifu/_0444_ ) );
INV_X1 \myifu/_1332_ ( .A(\myifu/_0177_ ), .ZN(\myifu/_0445_ ) );
OAI21_X1 \myifu/_1333_ ( .A(\myifu/_0443_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0445_ ), .ZN(\myifu/_0118_ ) );
OR2_X1 \myifu/_1334_ ( .A1(fanout_net_19 ), .A2(\myifu/_0146_ ), .ZN(\myifu/_0446_ ) );
AND3_X1 \myifu/_1335_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0901_ ), .ZN(\myifu/_0447_ ) );
OAI211_X2 \myifu/_1336_ ( .A(\myifu/_0437_ ), .B(\myifu/_0446_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0447_ ), .ZN(\myifu/_0448_ ) );
INV_X1 \myifu/_1337_ ( .A(\myifu/_0178_ ), .ZN(\myifu/_0449_ ) );
OAI21_X1 \myifu/_1338_ ( .A(\myifu/_0448_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0449_ ), .ZN(\myifu/_0119_ ) );
OAI21_X1 \myifu/_1339_ ( .A(\myifu/_0179_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0450_ ) );
OR2_X1 \myifu/_1340_ ( .A1(fanout_net_19 ), .A2(\myifu/_0147_ ), .ZN(\myifu/_0451_ ) );
AND3_X1 \myifu/_1341_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0902_ ), .ZN(\myifu/_0452_ ) );
OAI211_X2 \myifu/_1342_ ( .A(\myifu/_0428_ ), .B(\myifu/_0451_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0452_ ), .ZN(\myifu/_0453_ ) );
NAND2_X1 \myifu/_1343_ ( .A1(\myifu/_0450_ ), .A2(\myifu/_0453_ ), .ZN(\myifu/_0120_ ) );
OAI21_X1 \myifu/_1344_ ( .A(\myifu/_0180_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0454_ ) );
OR2_X1 \myifu/_1345_ ( .A1(fanout_net_19 ), .A2(\myifu/_0148_ ), .ZN(\myifu/_0455_ ) );
AND3_X1 \myifu/_1346_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0903_ ), .ZN(\myifu/_0456_ ) );
OAI211_X2 \myifu/_1347_ ( .A(\myifu/_0428_ ), .B(\myifu/_0455_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0456_ ), .ZN(\myifu/_0457_ ) );
NAND2_X1 \myifu/_1348_ ( .A1(\myifu/_0454_ ), .A2(\myifu/_0457_ ), .ZN(\myifu/_0121_ ) );
OR2_X1 \myifu/_1349_ ( .A1(fanout_net_19 ), .A2(\myifu/_0149_ ), .ZN(\myifu/_0458_ ) );
AND3_X1 \myifu/_1350_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0904_ ), .ZN(\myifu/_0459_ ) );
OAI211_X2 \myifu/_1351_ ( .A(\myifu/_0437_ ), .B(\myifu/_0458_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0459_ ), .ZN(\myifu/_0460_ ) );
INV_X1 \myifu/_1352_ ( .A(\myifu/_0181_ ), .ZN(\myifu/_0461_ ) );
OAI21_X1 \myifu/_1353_ ( .A(\myifu/_0460_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0461_ ), .ZN(\myifu/_0122_ ) );
OR2_X1 \myifu/_1354_ ( .A1(fanout_net_19 ), .A2(\myifu/_0150_ ), .ZN(\myifu/_0462_ ) );
AND3_X1 \myifu/_1355_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0905_ ), .ZN(\myifu/_0463_ ) );
OAI211_X2 \myifu/_1356_ ( .A(\myifu/_0437_ ), .B(\myifu/_0462_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0463_ ), .ZN(\myifu/_0464_ ) );
INV_X1 \myifu/_1357_ ( .A(\myifu/_0182_ ), .ZN(\myifu/_0465_ ) );
OAI21_X1 \myifu/_1358_ ( .A(\myifu/_0464_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0465_ ), .ZN(\myifu/_0123_ ) );
OR2_X1 \myifu/_1359_ ( .A1(fanout_net_19 ), .A2(\myifu/_0151_ ), .ZN(\myifu/_0466_ ) );
AND3_X1 \myifu/_1360_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0906_ ), .ZN(\myifu/_0467_ ) );
OAI211_X2 \myifu/_1361_ ( .A(\myifu/_0437_ ), .B(\myifu/_0466_ ), .C1(\myifu/_0358_ ), .C2(\myifu/_0467_ ), .ZN(\myifu/_0468_ ) );
INV_X1 \myifu/_1362_ ( .A(\myifu/_0183_ ), .ZN(\myifu/_0469_ ) );
OAI21_X1 \myifu/_1363_ ( .A(\myifu/_0468_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0469_ ), .ZN(\myifu/_0124_ ) );
OR2_X1 \myifu/_1364_ ( .A1(fanout_net_19 ), .A2(\myifu/_0152_ ), .ZN(\myifu/_0470_ ) );
AND3_X1 \myifu/_1365_ ( .A1(\myifu/_0351_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0907_ ), .ZN(\myifu/_0471_ ) );
OAI211_X2 \myifu/_1366_ ( .A(\myifu/_0437_ ), .B(\myifu/_0470_ ), .C1(\myifu/_0358_ ), .C2(\myifu/_0471_ ), .ZN(\myifu/_0472_ ) );
INV_X1 \myifu/_1367_ ( .A(\myifu/_0184_ ), .ZN(\myifu/_0473_ ) );
OAI21_X1 \myifu/_1368_ ( .A(\myifu/_0472_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0473_ ), .ZN(\myifu/_0125_ ) );
OAI21_X1 \myifu/_1369_ ( .A(\myifu/_0186_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0474_ ) );
OR2_X1 \myifu/_1370_ ( .A1(fanout_net_19 ), .A2(\myifu/_0154_ ), .ZN(\myifu/_0475_ ) );
AND3_X1 \myifu/_1371_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0909_ ), .ZN(\myifu/_0476_ ) );
OAI211_X2 \myifu/_1372_ ( .A(\myifu/_0428_ ), .B(\myifu/_0475_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0476_ ), .ZN(\myifu/_0477_ ) );
NAND2_X1 \myifu/_1373_ ( .A1(\myifu/_0474_ ), .A2(\myifu/_0477_ ), .ZN(\myifu/_0126_ ) );
OAI21_X1 \myifu/_1374_ ( .A(\myifu/_0187_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0478_ ) );
OR2_X1 \myifu/_1375_ ( .A1(fanout_net_19 ), .A2(\myifu/_0155_ ), .ZN(\myifu/_0479_ ) );
AND3_X1 \myifu/_1376_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0910_ ), .ZN(\myifu/_0480_ ) );
OAI211_X2 \myifu/_1377_ ( .A(\myifu/_0428_ ), .B(\myifu/_0479_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0480_ ), .ZN(\myifu/_0481_ ) );
NAND2_X1 \myifu/_1378_ ( .A1(\myifu/_0478_ ), .A2(\myifu/_0481_ ), .ZN(\myifu/_0127_ ) );
OR2_X1 \myifu/_1379_ ( .A1(fanout_net_19 ), .A2(\myifu/_0156_ ), .ZN(\myifu/_0482_ ) );
AND3_X1 \myifu/_1380_ ( .A1(\myifu/_0351_ ), .A2(\myifu/_0377_ ), .A3(\myifu/_0911_ ), .ZN(\myifu/_0483_ ) );
OAI211_X2 \myifu/_1381_ ( .A(\myifu/_0381_ ), .B(\myifu/_0482_ ), .C1(\myifu/_0358_ ), .C2(\myifu/_0483_ ), .ZN(\myifu/_0484_ ) );
INV_X1 \myifu/_1382_ ( .A(\myifu/_0188_ ), .ZN(\myifu/_0485_ ) );
OAI21_X1 \myifu/_1383_ ( .A(\myifu/_0484_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0485_ ), .ZN(\myifu/_0128_ ) );
OAI21_X1 \myifu/_1384_ ( .A(\myifu/_0189_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0486_ ) );
OR2_X1 \myifu/_1385_ ( .A1(fanout_net_19 ), .A2(\myifu/_0157_ ), .ZN(\myifu/_0487_ ) );
AND3_X1 \myifu/_1386_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0912_ ), .ZN(\myifu/_0488_ ) );
OAI211_X2 \myifu/_1387_ ( .A(\myifu/_0428_ ), .B(\myifu/_0487_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0488_ ), .ZN(\myifu/_0489_ ) );
NAND2_X1 \myifu/_1388_ ( .A1(\myifu/_0486_ ), .A2(\myifu/_0489_ ), .ZN(\myifu/_0129_ ) );
OAI21_X1 \myifu/_1389_ ( .A(\myifu/_0190_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0490_ ) );
OR2_X1 \myifu/_1390_ ( .A1(fanout_net_19 ), .A2(\myifu/_0158_ ), .ZN(\myifu/_0491_ ) );
AND3_X1 \myifu/_1391_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0913_ ), .ZN(\myifu/_0492_ ) );
OAI211_X2 \myifu/_1392_ ( .A(\myifu/_0428_ ), .B(\myifu/_0491_ ), .C1(\myifu/_0417_ ), .C2(\myifu/_0492_ ), .ZN(\myifu/_0493_ ) );
NAND2_X1 \myifu/_1393_ ( .A1(\myifu/_0490_ ), .A2(\myifu/_0493_ ), .ZN(\myifu/_0130_ ) );
OAI21_X1 \myifu/_1394_ ( .A(\myifu/_0191_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0494_ ) );
OR2_X1 \myifu/_1395_ ( .A1(fanout_net_19 ), .A2(\myifu/_0159_ ), .ZN(\myifu/_0495_ ) );
AND3_X1 \myifu/_1396_ ( .A1(\myifu/_0422_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0914_ ), .ZN(\myifu/_0496_ ) );
OAI211_X2 \myifu/_1397_ ( .A(\myifu/_0428_ ), .B(\myifu/_0495_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0496_ ), .ZN(\myifu/_0497_ ) );
NAND2_X1 \myifu/_1398_ ( .A1(\myifu/_0494_ ), .A2(\myifu/_0497_ ), .ZN(\myifu/_0131_ ) );
OAI21_X1 \myifu/_1399_ ( .A(\myifu/_0192_ ), .B1(\myifu/_0425_ ), .B2(\myifu/_0426_ ), .ZN(\myifu/_0498_ ) );
OR2_X1 \myifu/_1400_ ( .A1(fanout_net_19 ), .A2(\myifu/_0160_ ), .ZN(\myifu/_0499_ ) );
AND3_X1 \myifu/_1401_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0430_ ), .A3(\myifu/_0915_ ), .ZN(\myifu/_0500_ ) );
OAI211_X2 \myifu/_1402_ ( .A(\myifu/_0428_ ), .B(\myifu/_0499_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0500_ ), .ZN(\myifu/_0501_ ) );
NAND2_X1 \myifu/_1403_ ( .A1(\myifu/_0498_ ), .A2(\myifu/_0501_ ), .ZN(\myifu/_0132_ ) );
OAI21_X1 \myifu/_1404_ ( .A(\myifu/_0193_ ), .B1(\myifu/_0371_ ), .B2(\myifu/_0378_ ), .ZN(\myifu/_0502_ ) );
OR2_X1 \myifu/_1405_ ( .A1(\myifu/_0944_ ), .A2(\myifu/_0161_ ), .ZN(\myifu/_0503_ ) );
AND3_X1 \myifu/_1406_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0916_ ), .ZN(\myifu/_0504_ ) );
OAI211_X2 \myifu/_1407_ ( .A(\myifu/_0437_ ), .B(\myifu/_0503_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0504_ ), .ZN(\myifu/_0505_ ) );
NAND2_X1 \myifu/_1408_ ( .A1(\myifu/_0502_ ), .A2(\myifu/_0505_ ), .ZN(\myifu/_0133_ ) );
OAI21_X1 \myifu/_1409_ ( .A(\myifu/_0194_ ), .B1(\myifu/_0371_ ), .B2(\myifu/_0378_ ), .ZN(\myifu/_0506_ ) );
OR2_X1 \myifu/_1410_ ( .A1(\myifu/_0944_ ), .A2(\myifu/_0162_ ), .ZN(\myifu/_0507_ ) );
AND3_X1 \myifu/_1411_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0917_ ), .ZN(\myifu/_0508_ ) );
OAI211_X2 \myifu/_1412_ ( .A(\myifu/_0437_ ), .B(\myifu/_0507_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0508_ ), .ZN(\myifu/_0509_ ) );
NAND2_X1 \myifu/_1413_ ( .A1(\myifu/_0506_ ), .A2(\myifu/_0509_ ), .ZN(\myifu/_0134_ ) );
OAI21_X1 \myifu/_1414_ ( .A(\myifu/_0195_ ), .B1(\myifu/_0371_ ), .B2(\myifu/_0378_ ), .ZN(\myifu/_0510_ ) );
OR2_X1 \myifu/_1415_ ( .A1(\myifu/_0944_ ), .A2(\myifu/_0163_ ), .ZN(\myifu/_0511_ ) );
AND3_X1 \myifu/_1416_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0918_ ), .ZN(\myifu/_0512_ ) );
OAI211_X2 \myifu/_1417_ ( .A(\myifu/_0437_ ), .B(\myifu/_0511_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0512_ ), .ZN(\myifu/_0513_ ) );
NAND2_X1 \myifu/_1418_ ( .A1(\myifu/_0510_ ), .A2(\myifu/_0513_ ), .ZN(\myifu/_0135_ ) );
OAI21_X1 \myifu/_1419_ ( .A(\myifu/_0197_ ), .B1(\myifu/_0371_ ), .B2(\myifu/_0378_ ), .ZN(\myifu/_0514_ ) );
OR2_X1 \myifu/_1420_ ( .A1(\myifu/_0944_ ), .A2(\myifu/_0165_ ), .ZN(\myifu/_0515_ ) );
AND3_X1 \myifu/_1421_ ( .A1(\myifu/_0440_ ), .A2(\myifu/_0441_ ), .A3(\myifu/_0920_ ), .ZN(\myifu/_0516_ ) );
OAI211_X2 \myifu/_1422_ ( .A(\myifu/_0437_ ), .B(\myifu/_0515_ ), .C1(\myifu/_0439_ ), .C2(\myifu/_0516_ ), .ZN(\myifu/_0517_ ) );
NAND2_X1 \myifu/_1423_ ( .A1(\myifu/_0514_ ), .A2(\myifu/_0517_ ), .ZN(\myifu/_0136_ ) );
OR2_X1 \myifu/_1424_ ( .A1(\myifu/_0944_ ), .A2(\myifu/_0166_ ), .ZN(\myifu/_0518_ ) );
AND3_X1 \myifu/_1425_ ( .A1(\myifu/_0351_ ), .A2(\myifu/_0377_ ), .A3(\myifu/_0921_ ), .ZN(\myifu/_0519_ ) );
OAI211_X2 \myifu/_1426_ ( .A(\myifu/_0381_ ), .B(\myifu/_0518_ ), .C1(\myifu/_0358_ ), .C2(\myifu/_0519_ ), .ZN(\myifu/_0520_ ) );
INV_X32 \myifu/_1427_ ( .A(\myifu/_0896_ ), .ZN(\myifu/_0521_ ) );
OAI21_X1 \myifu/_1428_ ( .A(\myifu/_0520_ ), .B1(\myifu/_0444_ ), .B2(\myifu/_0521_ ), .ZN(\myifu/_0137_ ) );
MUX2_X1 \myifu/_1429_ ( .A(\myifu/_0365_ ), .B(\myifu/_0344_ ), .S(\myifu/_0943_ ), .Z(\myifu/_0522_ ) );
OAI21_X1 \myifu/_1430_ ( .A(\myifu/_0140_ ), .B1(\myifu/_0522_ ), .B2(fanout_net_18 ), .ZN(\myifu/_0523_ ) );
INV_X1 \myifu/_1431_ ( .A(\myifu/_0362_ ), .ZN(\myifu/_0524_ ) );
BUF_X4 \myifu/_1432_ ( .A(\myifu/_0524_ ), .Z(\myifu/_0525_ ) );
BUF_X4 \myifu/_1433_ ( .A(\myifu/_0525_ ), .Z(\myifu/_0526_ ) );
OAI21_X1 \myifu/_1434_ ( .A(\myifu/_0523_ ), .B1(fanout_net_18 ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0139_ ) );
AND2_X1 \myifu/_1435_ ( .A1(\myifu/_0281_ ), .A2(\myifu/_0141_ ), .ZN(\myifu/_0527_ ) );
INV_X1 \myifu/_1436_ ( .A(\myifu/_0527_ ), .ZN(\myifu/_0528_ ) );
NOR3_X1 \myifu/_1437_ ( .A1(\myifu/_0528_ ), .A2(\myifu/_0864_ ), .A3(\myifu/_0524_ ), .ZN(\myifu/_0529_ ) );
AND2_X1 \myifu/_1438_ ( .A1(\myifu/_0527_ ), .A2(\myifu/_0362_ ), .ZN(\myifu/_0530_ ) );
BUF_X4 \myifu/_1439_ ( .A(\myifu/_0530_ ), .Z(\myifu/_0531_ ) );
INV_X1 \myifu/_1440_ ( .A(\myifu/_0531_ ), .ZN(\myifu/_0532_ ) );
AOI211_X4 \myifu/_1441_ ( .A(fanout_net_18 ), .B(\myifu/_0529_ ), .C1(\myifu/_0366_ ), .C2(\myifu/_0532_ ), .ZN(\myifu/_0073_ ) );
NOR3_X4 \myifu/_1442_ ( .A1(\myifu/_0521_ ), .A2(\myifu/_0196_ ), .A3(\myifu/_0198_ ), .ZN(\myifu/_0533_ ) );
NAND3_X4 \myifu/_1443_ ( .A1(\myifu/_0533_ ), .A2(\myifu/_0174_ ), .A3(\myifu/_0185_ ), .ZN(\myifu/_0534_ ) );
NAND2_X4 \myifu/_1444_ ( .A1(\myifu/_0200_ ), .A2(\myifu/_0201_ ), .ZN(\myifu/_0535_ ) );
NOR2_X4 \myifu/_1445_ ( .A1(\myifu/_0535_ ), .A2(\myifu/_0199_ ), .ZN(\myifu/_0536_ ) );
INV_X4 \myifu/_1446_ ( .A(\myifu/_0536_ ), .ZN(\myifu/_0537_ ) );
NOR3_X1 \myifu/_1447_ ( .A1(\myifu/_0534_ ), .A2(\myifu/_0028_ ), .A3(\myifu/_0537_ ), .ZN(\myifu/_0538_ ) );
AND4_X4 \myifu/_1448_ ( .A1(\myifu/_0174_ ), .A2(\myifu/_0185_ ), .A3(\myifu/_0196_ ), .A4(\myifu/_0198_ ), .ZN(\myifu/_0539_ ) );
BUF_X8 \myifu/_1449_ ( .A(\myifu/_0536_ ), .Z(\myifu/_0540_ ) );
AND3_X1 \myifu/_1450_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0187_ ), .ZN(\myifu/_0541_ ) );
NOR2_X1 \myifu/_1451_ ( .A1(\myifu/_0538_ ), .A2(\myifu/_0541_ ), .ZN(\myifu/_0542_ ) );
XOR2_X1 \myifu/_1452_ ( .A(\myifu/_0542_ ), .B(\myifu/_0027_ ), .Z(\myifu/_0543_ ) );
AND2_X1 \myifu/_1453_ ( .A1(\myifu/_0528_ ), .A2(\myifu/_0543_ ), .ZN(\myifu/_0544_ ) );
AOI211_X4 \myifu/_1454_ ( .A(\myifu/_0524_ ), .B(\myifu/_0544_ ), .C1(\myifu/_0875_ ), .C2(\myifu/_0527_ ), .ZN(\myifu/_0545_ ) );
AOI211_X4 \myifu/_1455_ ( .A(fanout_net_18 ), .B(\myifu/_0545_ ), .C1(\myifu/_0367_ ), .C2(\myifu/_0525_ ), .ZN(\myifu/_0074_ ) );
OR2_X1 \myifu/_1456_ ( .A1(\myifu/_0528_ ), .A2(\myifu/_0886_ ), .ZN(\myifu/_0546_ ) );
BUF_X4 \myifu/_1457_ ( .A(\myifu/_0362_ ), .Z(\myifu/_0547_ ) );
BUF_X4 \myifu/_1458_ ( .A(\myifu/_0527_ ), .Z(\myifu/_0548_ ) );
NOR2_X4 \myifu/_1459_ ( .A1(\myifu/_0534_ ), .A2(\myifu/_0537_ ), .ZN(\myifu/_0549_ ) );
NAND2_X2 \myifu/_1460_ ( .A1(\myifu/_0549_ ), .A2(\myifu/_0029_ ), .ZN(\myifu/_0550_ ) );
NAND3_X1 \myifu/_1461_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0485_ ), .ZN(\myifu/_0551_ ) );
AND3_X4 \myifu/_1462_ ( .A1(\myifu/_0550_ ), .A2(\myifu/_0863_ ), .A3(\myifu/_0551_ ), .ZN(\myifu/_0552_ ) );
AOI21_X4 \myifu/_1463_ ( .A(\myifu/_0863_ ), .B1(\myifu/_0550_ ), .B2(\myifu/_0551_ ), .ZN(\myifu/_0553_ ) );
NOR2_X4 \myifu/_1464_ ( .A1(\myifu/_0552_ ), .A2(\myifu/_0553_ ), .ZN(\myifu/_0554_ ) );
NOR2_X1 \myifu/_1465_ ( .A1(\myifu/_0542_ ), .A2(\myifu/_0027_ ), .ZN(\myifu/_0555_ ) );
XOR2_X1 \myifu/_1466_ ( .A(\myifu/_0554_ ), .B(\myifu/_0555_ ), .Z(\myifu/_0556_ ) );
OAI211_X2 \myifu/_1467_ ( .A(\myifu/_0546_ ), .B(\myifu/_0547_ ), .C1(\myifu/_0548_ ), .C2(\myifu/_0556_ ), .ZN(\myifu/_0557_ ) );
OAI21_X1 \myifu/_1468_ ( .A(\myifu/_0863_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0558_ ) );
AOI21_X1 \myifu/_1469_ ( .A(fanout_net_18 ), .B1(\myifu/_0557_ ), .B2(\myifu/_0558_ ), .ZN(\myifu/_0075_ ) );
AND2_X1 \myifu/_1470_ ( .A1(\myifu/_0554_ ), .A2(\myifu/_0555_ ), .ZN(\myifu/_0559_ ) );
NAND3_X1 \myifu/_1471_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0189_ ), .ZN(\myifu/_0560_ ) );
INV_X4 \myifu/_1472_ ( .A(\myifu/_0549_ ), .ZN(\myifu/_0561_ ) );
BUF_X8 \myifu/_1473_ ( .A(\myifu/_0561_ ), .Z(\myifu/_0562_ ) );
OAI21_X2 \myifu/_1474_ ( .A(\myifu/_0560_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0030_ ), .ZN(\myifu/_0563_ ) );
XNOR2_X1 \myifu/_1475_ ( .A(\myifu/_0563_ ), .B(\myifu/_0266_ ), .ZN(\myifu/_0564_ ) );
OR3_X1 \myifu/_1476_ ( .A1(\myifu/_0559_ ), .A2(\myifu/_0552_ ), .A3(\myifu/_0564_ ), .ZN(\myifu/_0565_ ) );
OAI21_X1 \myifu/_1477_ ( .A(\myifu/_0564_ ), .B1(\myifu/_0559_ ), .B2(\myifu/_0552_ ), .ZN(\myifu/_0566_ ) );
NOR2_X2 \myifu/_1478_ ( .A1(\myifu/_0548_ ), .A2(\myifu/_0524_ ), .ZN(\myifu/_0567_ ) );
NAND3_X1 \myifu/_1479_ ( .A1(\myifu/_0565_ ), .A2(\myifu/_0566_ ), .A3(\myifu/_0567_ ), .ZN(\myifu/_0568_ ) );
BUF_X4 \myifu/_1480_ ( .A(\myifu/_0531_ ), .Z(\myifu/_0569_ ) );
AOI22_X1 \myifu/_1481_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0889_ ), .B1(\myifu/_0064_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0570_ ) );
AOI21_X1 \myifu/_1482_ ( .A(fanout_net_18 ), .B1(\myifu/_0568_ ), .B2(\myifu/_0570_ ), .ZN(\myifu/_0076_ ) );
BUF_X4 \myifu/_1483_ ( .A(\myifu/_0528_ ), .Z(\myifu/_0571_ ) );
AND2_X2 \myifu/_1484_ ( .A1(\myifu/_0563_ ), .A2(\myifu/_0064_ ), .ZN(\myifu/_0572_ ) );
INV_X1 \myifu/_1485_ ( .A(\myifu/_0572_ ), .ZN(\myifu/_0573_ ) );
NAND3_X1 \myifu/_1486_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0190_ ), .ZN(\myifu/_0574_ ) );
OAI21_X4 \myifu/_1487_ ( .A(\myifu/_0574_ ), .B1(\myifu/_0561_ ), .B2(\myifu/_0031_ ), .ZN(\myifu/_0575_ ) );
XOR2_X2 \myifu/_1488_ ( .A(\myifu/_0575_ ), .B(\myifu/_0065_ ), .Z(\myifu/_0576_ ) );
NAND3_X1 \myifu/_1489_ ( .A1(\myifu/_0566_ ), .A2(\myifu/_0573_ ), .A3(\myifu/_0576_ ), .ZN(\myifu/_0577_ ) );
NAND2_X1 \myifu/_1490_ ( .A1(\myifu/_0577_ ), .A2(\myifu/_0571_ ), .ZN(\myifu/_0578_ ) );
AOI21_X1 \myifu/_1491_ ( .A(\myifu/_0576_ ), .B1(\myifu/_0566_ ), .B2(\myifu/_0573_ ), .ZN(\myifu/_0579_ ) );
OAI221_X1 \myifu/_1492_ ( .A(\myifu/_0547_ ), .B1(\myifu/_0890_ ), .B2(\myifu/_0571_ ), .C1(\myifu/_0578_ ), .C2(\myifu/_0579_ ), .ZN(\myifu/_0580_ ) );
OAI21_X1 \myifu/_1493_ ( .A(\myifu/_0065_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0581_ ) );
AOI21_X1 \myifu/_1494_ ( .A(fanout_net_18 ), .B1(\myifu/_0580_ ), .B2(\myifu/_0581_ ), .ZN(\myifu/_0077_ ) );
AND2_X2 \myifu/_1495_ ( .A1(\myifu/_0576_ ), .A2(\myifu/_0572_ ), .ZN(\myifu/_0582_ ) );
AOI21_X1 \myifu/_1496_ ( .A(\myifu/_0582_ ), .B1(\myifu/_0065_ ), .B2(\myifu/_0575_ ), .ZN(\myifu/_0583_ ) );
OAI211_X2 \myifu/_1497_ ( .A(\myifu/_0564_ ), .B(\myifu/_0576_ ), .C1(\myifu/_0559_ ), .C2(\myifu/_0552_ ), .ZN(\myifu/_0584_ ) );
AND2_X4 \myifu/_1498_ ( .A1(\myifu/_0583_ ), .A2(\myifu/_0584_ ), .ZN(\myifu/_0585_ ) );
AND2_X4 \myifu/_1499_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .ZN(\myifu/_0586_ ) );
INV_X4 \myifu/_1500_ ( .A(\myifu/_0586_ ), .ZN(\myifu/_0587_ ) );
AOI21_X1 \myifu/_1501_ ( .A(\myifu/_0032_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0587_ ), .ZN(\myifu/_0588_ ) );
XNOR2_X1 \myifu/_1502_ ( .A(\myifu/_0588_ ), .B(\myifu/_0293_ ), .ZN(\myifu/_0589_ ) );
INV_X1 \myifu/_1503_ ( .A(\myifu/_0589_ ), .ZN(\myifu/_0590_ ) );
OR2_X1 \myifu/_1504_ ( .A1(\myifu/_0585_ ), .A2(\myifu/_0590_ ), .ZN(\myifu/_0591_ ) );
BUF_X4 \myifu/_1505_ ( .A(\myifu/_0567_ ), .Z(\myifu/_0592_ ) );
NAND3_X1 \myifu/_1506_ ( .A1(\myifu/_0583_ ), .A2(\myifu/_0584_ ), .A3(\myifu/_0590_ ), .ZN(\myifu/_0593_ ) );
NAND3_X1 \myifu/_1507_ ( .A1(\myifu/_0591_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0593_ ), .ZN(\myifu/_0594_ ) );
AOI22_X1 \myifu/_1508_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0891_ ), .B1(\myifu/_0066_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0595_ ) );
AOI21_X1 \myifu/_1509_ ( .A(fanout_net_18 ), .B1(\myifu/_0594_ ), .B2(\myifu/_0595_ ), .ZN(\myifu/_0078_ ) );
AND2_X2 \myifu/_1510_ ( .A1(\myifu/_0588_ ), .A2(\myifu/_0066_ ), .ZN(\myifu/_0596_ ) );
INV_X1 \myifu/_1511_ ( .A(\myifu/_0596_ ), .ZN(\myifu/_0597_ ) );
AOI21_X2 \myifu/_1512_ ( .A(\myifu/_0033_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0587_ ), .ZN(\myifu/_0598_ ) );
NOR2_X1 \myifu/_1513_ ( .A1(\myifu/_0598_ ), .A2(\myifu/_0067_ ), .ZN(\myifu/_0599_ ) );
NOR2_X4 \myifu/_1514_ ( .A1(\myifu/_0549_ ), .A2(\myifu/_0586_ ), .ZN(\myifu/_0600_ ) );
NOR3_X4 \myifu/_1515_ ( .A1(\myifu/_0600_ ), .A2(\myifu/_0282_ ), .A3(\myifu/_0033_ ), .ZN(\myifu/_0601_ ) );
NOR2_X4 \myifu/_1516_ ( .A1(\myifu/_0599_ ), .A2(\myifu/_0601_ ), .ZN(\myifu/_0602_ ) );
NAND3_X1 \myifu/_1517_ ( .A1(\myifu/_0591_ ), .A2(\myifu/_0597_ ), .A3(\myifu/_0602_ ), .ZN(\myifu/_0603_ ) );
NAND2_X1 \myifu/_1518_ ( .A1(\myifu/_0603_ ), .A2(\myifu/_0571_ ), .ZN(\myifu/_0604_ ) );
AOI21_X1 \myifu/_1519_ ( .A(\myifu/_0602_ ), .B1(\myifu/_0591_ ), .B2(\myifu/_0597_ ), .ZN(\myifu/_0605_ ) );
OAI221_X1 \myifu/_1520_ ( .A(\myifu/_0547_ ), .B1(\myifu/_0892_ ), .B2(\myifu/_0571_ ), .C1(\myifu/_0604_ ), .C2(\myifu/_0605_ ), .ZN(\myifu/_0606_ ) );
OAI21_X1 \myifu/_1521_ ( .A(\myifu/_0067_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0607_ ) );
AOI21_X1 \myifu/_1522_ ( .A(fanout_net_18 ), .B1(\myifu/_0606_ ), .B2(\myifu/_0607_ ), .ZN(\myifu/_0079_ ) );
NOR4_X1 \myifu/_1523_ ( .A1(\myifu/_0585_ ), .A2(\myifu/_0590_ ), .A3(\myifu/_0601_ ), .A4(\myifu/_0599_ ), .ZN(\myifu/_0608_ ) );
AOI21_X4 \myifu/_1524_ ( .A(\myifu/_0034_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0587_ ), .ZN(\myifu/_0609_ ) );
XOR2_X2 \myifu/_1525_ ( .A(\myifu/_0609_ ), .B(\myifu/_0068_ ), .Z(\myifu/_0610_ ) );
AOI21_X1 \myifu/_1526_ ( .A(\myifu/_0601_ ), .B1(\myifu/_0602_ ), .B2(\myifu/_0596_ ), .ZN(\myifu/_0611_ ) );
INV_X2 \myifu/_1527_ ( .A(\myifu/_0611_ ), .ZN(\myifu/_0612_ ) );
OR3_X1 \myifu/_1528_ ( .A1(\myifu/_0608_ ), .A2(\myifu/_0610_ ), .A3(\myifu/_0612_ ), .ZN(\myifu/_0613_ ) );
OAI21_X1 \myifu/_1529_ ( .A(\myifu/_0610_ ), .B1(\myifu/_0608_ ), .B2(\myifu/_0612_ ), .ZN(\myifu/_0614_ ) );
NAND3_X1 \myifu/_1530_ ( .A1(\myifu/_0613_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0614_ ), .ZN(\myifu/_0615_ ) );
AOI22_X1 \myifu/_1531_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0893_ ), .B1(\myifu/_0068_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0616_ ) );
AOI21_X1 \myifu/_1532_ ( .A(fanout_net_18 ), .B1(\myifu/_0615_ ), .B2(\myifu/_0616_ ), .ZN(\myifu/_0080_ ) );
NAND2_X1 \myifu/_1533_ ( .A1(\myifu/_0609_ ), .A2(\myifu/_0068_ ), .ZN(\myifu/_0617_ ) );
NAND2_X1 \myifu/_1534_ ( .A1(\myifu/_0614_ ), .A2(\myifu/_0617_ ), .ZN(\myifu/_0618_ ) );
NOR3_X1 \myifu/_1535_ ( .A1(\myifu/_0600_ ), .A2(\myifu/_0305_ ), .A3(\myifu/_0035_ ), .ZN(\myifu/_0619_ ) );
INV_X1 \myifu/_1536_ ( .A(\myifu/_0619_ ), .ZN(\myifu/_0620_ ) );
OAI21_X1 \myifu/_1537_ ( .A(\myifu/_0305_ ), .B1(\myifu/_0600_ ), .B2(\myifu/_0035_ ), .ZN(\myifu/_0621_ ) );
AND2_X1 \myifu/_1538_ ( .A1(\myifu/_0620_ ), .A2(\myifu/_0621_ ), .ZN(\myifu/_0622_ ) );
INV_X1 \myifu/_1539_ ( .A(\myifu/_0622_ ), .ZN(\myifu/_0623_ ) );
OAI21_X1 \myifu/_1540_ ( .A(\myifu/_0571_ ), .B1(\myifu/_0618_ ), .B2(\myifu/_0623_ ), .ZN(\myifu/_0624_ ) );
AOI21_X1 \myifu/_1541_ ( .A(\myifu/_0622_ ), .B1(\myifu/_0614_ ), .B2(\myifu/_0617_ ), .ZN(\myifu/_0625_ ) );
OAI221_X1 \myifu/_1542_ ( .A(\myifu/_0547_ ), .B1(\myifu/_0894_ ), .B2(\myifu/_0571_ ), .C1(\myifu/_0624_ ), .C2(\myifu/_0625_ ), .ZN(\myifu/_0626_ ) );
OAI21_X1 \myifu/_1543_ ( .A(\myifu/_0069_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0627_ ) );
AOI21_X1 \myifu/_1544_ ( .A(fanout_net_18 ), .B1(\myifu/_0626_ ), .B2(\myifu/_0627_ ), .ZN(\myifu/_0081_ ) );
NAND4_X1 \myifu/_1545_ ( .A1(\myifu/_0610_ ), .A2(\myifu/_0622_ ), .A3(\myifu/_0589_ ), .A4(\myifu/_0602_ ), .ZN(\myifu/_0628_ ) );
OR2_X4 \myifu/_1546_ ( .A1(\myifu/_0585_ ), .A2(\myifu/_0628_ ), .ZN(\myifu/_0629_ ) );
NAND3_X1 \myifu/_1547_ ( .A1(\myifu/_0612_ ), .A2(\myifu/_0610_ ), .A3(\myifu/_0622_ ), .ZN(\myifu/_0630_ ) );
NAND4_X1 \myifu/_1548_ ( .A1(\myifu/_0620_ ), .A2(\myifu/_0068_ ), .A3(\myifu/_0609_ ), .A4(\myifu/_0621_ ), .ZN(\myifu/_0631_ ) );
AND3_X4 \myifu/_1549_ ( .A1(\myifu/_0630_ ), .A2(\myifu/_0620_ ), .A3(\myifu/_0631_ ), .ZN(\myifu/_0632_ ) );
AND2_X4 \myifu/_1550_ ( .A1(\myifu/_0629_ ), .A2(\myifu/_0632_ ), .ZN(\myifu/_0633_ ) );
AOI21_X1 \myifu/_1551_ ( .A(\myifu/_0036_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0587_ ), .ZN(\myifu/_0634_ ) );
INV_X1 \myifu/_1552_ ( .A(\myifu/_0070_ ), .ZN(\myifu/_0635_ ) );
XNOR2_X1 \myifu/_1553_ ( .A(\myifu/_0634_ ), .B(\myifu/_0635_ ), .ZN(\myifu/_0636_ ) );
INV_X1 \myifu/_1554_ ( .A(\myifu/_0636_ ), .ZN(\myifu/_0637_ ) );
NOR2_X1 \myifu/_1555_ ( .A1(\myifu/_0633_ ), .A2(\myifu/_0637_ ), .ZN(\myifu/_0638_ ) );
INV_X1 \myifu/_1556_ ( .A(\myifu/_0638_ ), .ZN(\myifu/_0639_ ) );
NAND3_X1 \myifu/_1557_ ( .A1(\myifu/_0629_ ), .A2(\myifu/_0632_ ), .A3(\myifu/_0637_ ), .ZN(\myifu/_0640_ ) );
NAND3_X1 \myifu/_1558_ ( .A1(\myifu/_0639_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0640_ ), .ZN(\myifu/_0641_ ) );
AOI22_X1 \myifu/_1559_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0895_ ), .B1(\myifu/_0070_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0642_ ) );
AOI21_X1 \myifu/_1560_ ( .A(fanout_net_18 ), .B1(\myifu/_0641_ ), .B2(\myifu/_0642_ ), .ZN(\myifu/_0082_ ) );
AND2_X1 \myifu/_1561_ ( .A1(\myifu/_0634_ ), .A2(\myifu/_0070_ ), .ZN(\myifu/_0643_ ) );
OR2_X1 \myifu/_1562_ ( .A1(\myifu/_0638_ ), .A2(\myifu/_0643_ ), .ZN(\myifu/_0644_ ) );
AOI21_X1 \myifu/_1563_ ( .A(\myifu/_0037_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0587_ ), .ZN(\myifu/_0645_ ) );
NOR2_X1 \myifu/_1564_ ( .A1(\myifu/_0645_ ), .A2(\myifu/_0042_ ), .ZN(\myifu/_0646_ ) );
NOR3_X1 \myifu/_1565_ ( .A1(\myifu/_0600_ ), .A2(\myifu/_0338_ ), .A3(\myifu/_0037_ ), .ZN(\myifu/_0647_ ) );
NOR2_X1 \myifu/_1566_ ( .A1(\myifu/_0646_ ), .A2(\myifu/_0647_ ), .ZN(\myifu/_0648_ ) );
INV_X1 \myifu/_1567_ ( .A(\myifu/_0648_ ), .ZN(\myifu/_0649_ ) );
AND2_X1 \myifu/_1568_ ( .A1(\myifu/_0644_ ), .A2(\myifu/_0649_ ), .ZN(\myifu/_0650_ ) );
OAI21_X1 \myifu/_1569_ ( .A(\myifu/_0528_ ), .B1(\myifu/_0644_ ), .B2(\myifu/_0649_ ), .ZN(\myifu/_0651_ ) );
OAI221_X1 \myifu/_1570_ ( .A(\myifu/_0547_ ), .B1(\myifu/_0865_ ), .B2(\myifu/_0571_ ), .C1(\myifu/_0650_ ), .C2(\myifu/_0651_ ), .ZN(\myifu/_0652_ ) );
OAI21_X1 \myifu/_1571_ ( .A(\myifu/_0042_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0653_ ) );
AOI21_X1 \myifu/_1572_ ( .A(fanout_net_18 ), .B1(\myifu/_0652_ ), .B2(\myifu/_0653_ ), .ZN(\myifu/_0083_ ) );
AOI21_X1 \myifu/_1573_ ( .A(\myifu/_0647_ ), .B1(\myifu/_0070_ ), .B2(\myifu/_0634_ ), .ZN(\myifu/_0654_ ) );
INV_X1 \myifu/_1574_ ( .A(\myifu/_0654_ ), .ZN(\myifu/_0655_ ) );
INV_X8 \myifu/_1575_ ( .A(\myifu/_0633_ ), .ZN(\myifu/_0656_ ) );
AOI21_X1 \myifu/_1576_ ( .A(\myifu/_0655_ ), .B1(\myifu/_0656_ ), .B2(\myifu/_0636_ ), .ZN(\myifu/_0657_ ) );
NAND3_X1 \myifu/_1577_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0186_ ), .ZN(\myifu/_0658_ ) );
OAI21_X4 \myifu/_1578_ ( .A(\myifu/_0658_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0038_ ), .ZN(\myifu/_0659_ ) );
XNOR2_X2 \myifu/_1579_ ( .A(\myifu/_0659_ ), .B(\myifu/_0298_ ), .ZN(\myifu/_0660_ ) );
INV_X1 \myifu/_1580_ ( .A(\myifu/_0660_ ), .ZN(\myifu/_0661_ ) );
OR3_X1 \myifu/_1581_ ( .A1(\myifu/_0657_ ), .A2(\myifu/_0646_ ), .A3(\myifu/_0661_ ), .ZN(\myifu/_0662_ ) );
OAI21_X1 \myifu/_1582_ ( .A(\myifu/_0661_ ), .B1(\myifu/_0657_ ), .B2(\myifu/_0646_ ), .ZN(\myifu/_0663_ ) );
NAND3_X1 \myifu/_1583_ ( .A1(\myifu/_0662_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0663_ ), .ZN(\myifu/_0664_ ) );
AOI22_X1 \myifu/_1584_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0866_ ), .B1(\myifu/_0043_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0665_ ) );
AOI21_X1 \myifu/_1585_ ( .A(fanout_net_18 ), .B1(\myifu/_0664_ ), .B2(\myifu/_0665_ ), .ZN(\myifu/_0084_ ) );
AND2_X1 \myifu/_1586_ ( .A1(\myifu/_0659_ ), .A2(\myifu/_0043_ ), .ZN(\myifu/_0666_ ) );
INV_X1 \myifu/_1587_ ( .A(\myifu/_0666_ ), .ZN(\myifu/_0667_ ) );
AND2_X1 \myifu/_1588_ ( .A1(\myifu/_0662_ ), .A2(\myifu/_0667_ ), .ZN(\myifu/_0668_ ) );
OAI22_X1 \myifu/_1589_ ( .A1(\myifu/_0587_ ), .A2(\myifu/_0445_ ), .B1(\myifu/_0537_ ), .B2(\myifu/_0534_ ), .ZN(\myifu/_0669_ ) );
NAND2_X4 \myifu/_1590_ ( .A1(\myifu/_0549_ ), .A2(\myifu/_0039_ ), .ZN(\myifu/_0670_ ) );
AND3_X1 \myifu/_1591_ ( .A1(\myifu/_0669_ ), .A2(\myifu/_0044_ ), .A3(\myifu/_0670_ ), .ZN(\myifu/_0671_ ) );
AOI21_X1 \myifu/_1592_ ( .A(\myifu/_0044_ ), .B1(\myifu/_0669_ ), .B2(\myifu/_0670_ ), .ZN(\myifu/_0672_ ) );
NOR2_X2 \myifu/_1593_ ( .A1(\myifu/_0671_ ), .A2(\myifu/_0672_ ), .ZN(\myifu/_0673_ ) );
XNOR2_X1 \myifu/_1594_ ( .A(\myifu/_0668_ ), .B(\myifu/_0673_ ), .ZN(\myifu/_0674_ ) );
AND3_X1 \myifu/_1595_ ( .A1(\myifu/_0867_ ), .A2(\myifu/_0943_ ), .A3(\myifu/_0929_ ), .ZN(\myifu/_0675_ ) );
OAI22_X1 \myifu/_1596_ ( .A1(\myifu/_0674_ ), .A2(\myifu/_0548_ ), .B1(\myifu/_0567_ ), .B2(\myifu/_0675_ ), .ZN(\myifu/_0676_ ) );
OAI21_X1 \myifu/_1597_ ( .A(\myifu/_0044_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0677_ ) );
AOI21_X1 \myifu/_1598_ ( .A(fanout_net_18 ), .B1(\myifu/_0676_ ), .B2(\myifu/_0677_ ), .ZN(\myifu/_0085_ ) );
AND2_X1 \myifu/_1599_ ( .A1(\myifu/_0636_ ), .A2(\myifu/_0648_ ), .ZN(\myifu/_0678_ ) );
AND2_X1 \myifu/_1600_ ( .A1(\myifu/_0660_ ), .A2(\myifu/_0673_ ), .ZN(\myifu/_0679_ ) );
AND3_X1 \myifu/_1601_ ( .A1(\myifu/_0656_ ), .A2(\myifu/_0678_ ), .A3(\myifu/_0679_ ), .ZN(\myifu/_0680_ ) );
OAI211_X2 \myifu/_1602_ ( .A(\myifu/_0660_ ), .B(\myifu/_0673_ ), .C1(\myifu/_0643_ ), .C2(\myifu/_0647_ ), .ZN(\myifu/_0681_ ) );
NOR2_X2 \myifu/_1603_ ( .A1(\myifu/_0681_ ), .A2(\myifu/_0646_ ), .ZN(\myifu/_0682_ ) );
AND2_X1 \myifu/_1604_ ( .A1(\myifu/_0673_ ), .A2(\myifu/_0666_ ), .ZN(\myifu/_0683_ ) );
NOR3_X2 \myifu/_1605_ ( .A1(\myifu/_0682_ ), .A2(\myifu/_0671_ ), .A3(\myifu/_0683_ ), .ZN(\myifu/_0684_ ) );
INV_X2 \myifu/_1606_ ( .A(\myifu/_0684_ ), .ZN(\myifu/_0685_ ) );
NOR2_X1 \myifu/_1607_ ( .A1(\myifu/_0680_ ), .A2(\myifu/_0685_ ), .ZN(\myifu/_0686_ ) );
AND2_X1 \myifu/_1608_ ( .A1(\myifu/_0549_ ), .A2(\myifu/_0039_ ), .ZN(\myifu/_0687_ ) );
NAND3_X1 \myifu/_1609_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0178_ ), .ZN(\myifu/_0688_ ) );
AOI21_X1 \myifu/_1610_ ( .A(\myifu/_0687_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0688_ ), .ZN(\myifu/_0689_ ) );
INV_X1 \myifu/_1611_ ( .A(\myifu/_0045_ ), .ZN(\myifu/_0690_ ) );
XNOR2_X1 \myifu/_1612_ ( .A(\myifu/_0689_ ), .B(\myifu/_0690_ ), .ZN(\myifu/_0691_ ) );
INV_X1 \myifu/_1613_ ( .A(\myifu/_0691_ ), .ZN(\myifu/_0692_ ) );
NOR2_X1 \myifu/_1614_ ( .A1(\myifu/_0686_ ), .A2(\myifu/_0692_ ), .ZN(\myifu/_0693_ ) );
INV_X1 \myifu/_1615_ ( .A(\myifu/_0693_ ), .ZN(\myifu/_0694_ ) );
OR3_X1 \myifu/_1616_ ( .A1(\myifu/_0680_ ), .A2(\myifu/_0685_ ), .A3(\myifu/_0691_ ), .ZN(\myifu/_0695_ ) );
NAND3_X1 \myifu/_1617_ ( .A1(\myifu/_0694_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0695_ ), .ZN(\myifu/_0696_ ) );
AOI22_X1 \myifu/_1618_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0868_ ), .B1(\myifu/_0045_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0697_ ) );
AOI21_X1 \myifu/_1619_ ( .A(fanout_net_18 ), .B1(\myifu/_0696_ ), .B2(\myifu/_0697_ ), .ZN(\myifu/_0086_ ) );
AND2_X1 \myifu/_1620_ ( .A1(\myifu/_0689_ ), .A2(\myifu/_0045_ ), .ZN(\myifu/_0698_ ) );
NOR2_X1 \myifu/_1621_ ( .A1(\myifu/_0693_ ), .A2(\myifu/_0698_ ), .ZN(\myifu/_0699_ ) );
AND3_X1 \myifu/_1622_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0179_ ), .ZN(\myifu/_0700_ ) );
OAI21_X2 \myifu/_1623_ ( .A(\myifu/_0670_ ), .B1(\myifu/_0549_ ), .B2(\myifu/_0700_ ), .ZN(\myifu/_0701_ ) );
XNOR2_X2 \myifu/_1624_ ( .A(\myifu/_0701_ ), .B(\myifu/_0046_ ), .ZN(\myifu/_0702_ ) );
XNOR2_X1 \myifu/_1625_ ( .A(\myifu/_0699_ ), .B(\myifu/_0702_ ), .ZN(\myifu/_0703_ ) );
NAND2_X1 \myifu/_1626_ ( .A1(\myifu/_0703_ ), .A2(\myifu/_0592_ ), .ZN(\myifu/_0704_ ) );
AOI22_X1 \myifu/_1627_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0869_ ), .B1(\myifu/_0046_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0705_ ) );
AOI21_X1 \myifu/_1628_ ( .A(fanout_net_18 ), .B1(\myifu/_0704_ ), .B2(\myifu/_0705_ ), .ZN(\myifu/_0087_ ) );
AOI21_X1 \myifu/_1629_ ( .A(\myifu/_0699_ ), .B1(\myifu/_0284_ ), .B2(\myifu/_0701_ ), .ZN(\myifu/_0706_ ) );
NOR2_X1 \myifu/_1630_ ( .A1(\myifu/_0701_ ), .A2(\myifu/_0284_ ), .ZN(\myifu/_0707_ ) );
AND3_X1 \myifu/_1631_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0180_ ), .ZN(\myifu/_0708_ ) );
OAI21_X2 \myifu/_1632_ ( .A(\myifu/_0670_ ), .B1(\myifu/_0549_ ), .B2(\myifu/_0708_ ), .ZN(\myifu/_0709_ ) );
XNOR2_X1 \myifu/_1633_ ( .A(\myifu/_0709_ ), .B(\myifu/_0047_ ), .ZN(\myifu/_0710_ ) );
OR3_X1 \myifu/_1634_ ( .A1(\myifu/_0706_ ), .A2(\myifu/_0707_ ), .A3(\myifu/_0710_ ), .ZN(\myifu/_0711_ ) );
OAI21_X1 \myifu/_1635_ ( .A(\myifu/_0710_ ), .B1(\myifu/_0706_ ), .B2(\myifu/_0707_ ), .ZN(\myifu/_0712_ ) );
NAND3_X1 \myifu/_1636_ ( .A1(\myifu/_0711_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0712_ ), .ZN(\myifu/_0713_ ) );
AOI22_X1 \myifu/_1637_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0870_ ), .B1(\myifu/_0047_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0714_ ) );
AOI21_X1 \myifu/_1638_ ( .A(fanout_net_18 ), .B1(\myifu/_0713_ ), .B2(\myifu/_0714_ ), .ZN(\myifu/_0088_ ) );
OR2_X1 \myifu/_1639_ ( .A1(\myifu/_0709_ ), .A2(\myifu/_0300_ ), .ZN(\myifu/_0715_ ) );
AND2_X1 \myifu/_1640_ ( .A1(\myifu/_0712_ ), .A2(\myifu/_0715_ ), .ZN(\myifu/_0716_ ) );
OAI22_X1 \myifu/_1641_ ( .A1(\myifu/_0587_ ), .A2(\myifu/_0461_ ), .B1(\myifu/_0537_ ), .B2(\myifu/_0534_ ), .ZN(\myifu/_0717_ ) );
AND3_X4 \myifu/_1642_ ( .A1(\myifu/_0717_ ), .A2(\myifu/_0048_ ), .A3(\myifu/_0670_ ), .ZN(\myifu/_0718_ ) );
AOI21_X1 \myifu/_1643_ ( .A(\myifu/_0048_ ), .B1(\myifu/_0717_ ), .B2(\myifu/_0670_ ), .ZN(\myifu/_0719_ ) );
NOR2_X1 \myifu/_1644_ ( .A1(\myifu/_0718_ ), .A2(\myifu/_0719_ ), .ZN(\myifu/_0720_ ) );
XNOR2_X1 \myifu/_1645_ ( .A(\myifu/_0716_ ), .B(\myifu/_0720_ ), .ZN(\myifu/_0721_ ) );
AND3_X1 \myifu/_1646_ ( .A1(\myifu/_0871_ ), .A2(\myifu/_0943_ ), .A3(\myifu/_0929_ ), .ZN(\myifu/_0722_ ) );
OAI22_X1 \myifu/_1647_ ( .A1(\myifu/_0721_ ), .A2(\myifu/_0548_ ), .B1(\myifu/_0567_ ), .B2(\myifu/_0722_ ), .ZN(\myifu/_0723_ ) );
OAI21_X1 \myifu/_1648_ ( .A(\myifu/_0048_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0724_ ) );
AOI21_X1 \myifu/_1649_ ( .A(fanout_net_18 ), .B1(\myifu/_0723_ ), .B2(\myifu/_0724_ ), .ZN(\myifu/_0089_ ) );
OAI22_X1 \myifu/_1650_ ( .A1(\myifu/_0587_ ), .A2(\myifu/_0465_ ), .B1(\myifu/_0537_ ), .B2(\myifu/_0534_ ), .ZN(\myifu/_0725_ ) );
NAND2_X1 \myifu/_1651_ ( .A1(\myifu/_0725_ ), .A2(\myifu/_0670_ ), .ZN(\myifu/_0726_ ) );
XNOR2_X1 \myifu/_1652_ ( .A(\myifu/_0726_ ), .B(\myifu/_0049_ ), .ZN(\myifu/_0727_ ) );
INV_X1 \myifu/_1653_ ( .A(\myifu/_0727_ ), .ZN(\myifu/_0728_ ) );
AND2_X1 \myifu/_1654_ ( .A1(\myifu/_0710_ ), .A2(\myifu/_0720_ ), .ZN(\myifu/_0729_ ) );
AND3_X4 \myifu/_1655_ ( .A1(\myifu/_0729_ ), .A2(\myifu/_0691_ ), .A3(\myifu/_0702_ ), .ZN(\myifu/_0730_ ) );
NAND4_X4 \myifu/_1656_ ( .A1(\myifu/_0656_ ), .A2(\myifu/_0678_ ), .A3(\myifu/_0679_ ), .A4(\myifu/_0730_ ), .ZN(\myifu/_0731_ ) );
AND2_X2 \myifu/_1657_ ( .A1(\myifu/_0685_ ), .A2(\myifu/_0730_ ), .ZN(\myifu/_0732_ ) );
NOR4_X1 \myifu/_1658_ ( .A1(\myifu/_0718_ ), .A2(\myifu/_0719_ ), .A3(\myifu/_0300_ ), .A4(\myifu/_0709_ ), .ZN(\myifu/_0733_ ) );
NAND2_X1 \myifu/_1659_ ( .A1(\myifu/_0702_ ), .A2(\myifu/_0698_ ), .ZN(\myifu/_0734_ ) );
OAI21_X1 \myifu/_1660_ ( .A(\myifu/_0734_ ), .B1(\myifu/_0284_ ), .B2(\myifu/_0701_ ), .ZN(\myifu/_0735_ ) );
AND2_X2 \myifu/_1661_ ( .A1(\myifu/_0735_ ), .A2(\myifu/_0729_ ), .ZN(\myifu/_0736_ ) );
NOR4_X4 \myifu/_1662_ ( .A1(\myifu/_0732_ ), .A2(\myifu/_0718_ ), .A3(\myifu/_0733_ ), .A4(\myifu/_0736_ ), .ZN(\myifu/_0737_ ) );
AOI21_X1 \myifu/_1663_ ( .A(\myifu/_0728_ ), .B1(\myifu/_0731_ ), .B2(\myifu/_0737_ ), .ZN(\myifu/_0738_ ) );
INV_X1 \myifu/_1664_ ( .A(\myifu/_0738_ ), .ZN(\myifu/_0739_ ) );
NAND3_X1 \myifu/_1665_ ( .A1(\myifu/_0731_ ), .A2(\myifu/_0737_ ), .A3(\myifu/_0728_ ), .ZN(\myifu/_0740_ ) );
NAND3_X1 \myifu/_1666_ ( .A1(\myifu/_0739_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0740_ ), .ZN(\myifu/_0741_ ) );
AOI22_X1 \myifu/_1667_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0872_ ), .B1(\myifu/_0049_ ), .B2(\myifu/_0526_ ), .ZN(\myifu/_0742_ ) );
AOI21_X1 \myifu/_1668_ ( .A(fanout_net_18 ), .B1(\myifu/_0741_ ), .B2(\myifu/_0742_ ), .ZN(\myifu/_0090_ ) );
OAI22_X1 \myifu/_1669_ ( .A1(\myifu/_0587_ ), .A2(\myifu/_0469_ ), .B1(\myifu/_0537_ ), .B2(\myifu/_0534_ ), .ZN(\myifu/_0743_ ) );
AND2_X1 \myifu/_1670_ ( .A1(\myifu/_0743_ ), .A2(\myifu/_0670_ ), .ZN(\myifu/_0744_ ) );
XNOR2_X1 \myifu/_1671_ ( .A(\myifu/_0744_ ), .B(\myifu/_0040_ ), .ZN(\myifu/_0745_ ) );
INV_X1 \myifu/_1672_ ( .A(\myifu/_0745_ ), .ZN(\myifu/_0746_ ) );
AND3_X1 \myifu/_1673_ ( .A1(\myifu/_0725_ ), .A2(\myifu/_0049_ ), .A3(\myifu/_0670_ ), .ZN(\myifu/_0747_ ) );
INV_X1 \myifu/_1674_ ( .A(\myifu/_0747_ ), .ZN(\myifu/_0748_ ) );
AOI21_X1 \myifu/_1675_ ( .A(\myifu/_0746_ ), .B1(\myifu/_0739_ ), .B2(\myifu/_0748_ ), .ZN(\myifu/_0749_ ) );
INV_X1 \myifu/_1676_ ( .A(\myifu/_0749_ ), .ZN(\myifu/_0750_ ) );
NAND3_X1 \myifu/_1677_ ( .A1(\myifu/_0739_ ), .A2(\myifu/_0748_ ), .A3(\myifu/_0746_ ), .ZN(\myifu/_0751_ ) );
NAND3_X1 \myifu/_1678_ ( .A1(\myifu/_0750_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0751_ ), .ZN(\myifu/_0752_ ) );
AOI22_X1 \myifu/_1679_ ( .A1(\myifu/_0569_ ), .A2(\myifu/_0873_ ), .B1(\myifu/_0050_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0753_ ) );
AOI21_X1 \myifu/_1680_ ( .A(fanout_net_18 ), .B1(\myifu/_0752_ ), .B2(\myifu/_0753_ ), .ZN(\myifu/_0091_ ) );
AND3_X1 \myifu/_1681_ ( .A1(\myifu/_0743_ ), .A2(\myifu/_0050_ ), .A3(\myifu/_0670_ ), .ZN(\myifu/_0754_ ) );
NAND3_X1 \myifu/_1682_ ( .A1(\myifu/_0539_ ), .A2(\myifu/_0540_ ), .A3(\myifu/_0184_ ), .ZN(\myifu/_0755_ ) );
AOI21_X2 \myifu/_1683_ ( .A(\myifu/_0687_ ), .B1(\myifu/_0562_ ), .B2(\myifu/_0755_ ), .ZN(\myifu/_0756_ ) );
XOR2_X1 \myifu/_1684_ ( .A(\myifu/_0756_ ), .B(\myifu/_0051_ ), .Z(\myifu/_0757_ ) );
OR3_X1 \myifu/_1685_ ( .A1(\myifu/_0749_ ), .A2(\myifu/_0754_ ), .A3(\myifu/_0757_ ), .ZN(\myifu/_0758_ ) );
OAI21_X1 \myifu/_1686_ ( .A(\myifu/_0757_ ), .B1(\myifu/_0749_ ), .B2(\myifu/_0754_ ), .ZN(\myifu/_0759_ ) );
NAND3_X1 \myifu/_1687_ ( .A1(\myifu/_0758_ ), .A2(\myifu/_0592_ ), .A3(\myifu/_0759_ ), .ZN(\myifu/_0760_ ) );
AOI22_X1 \myifu/_1688_ ( .A1(\myifu/_0531_ ), .A2(\myifu/_0874_ ), .B1(\myifu/_0051_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0761_ ) );
AOI21_X1 \myifu/_1689_ ( .A(fanout_net_18 ), .B1(\myifu/_0760_ ), .B2(\myifu/_0761_ ), .ZN(\myifu/_0092_ ) );
NAND2_X1 \myifu/_1690_ ( .A1(\myifu/_0756_ ), .A2(\myifu/_0051_ ), .ZN(\myifu/_0762_ ) );
AND2_X1 \myifu/_1691_ ( .A1(\myifu/_0759_ ), .A2(\myifu/_0762_ ), .ZN(\myifu/_0763_ ) );
NOR2_X2 \myifu/_1692_ ( .A1(\myifu/_0600_ ), .A2(\myifu/_0039_ ), .ZN(\myifu/_0764_ ) );
XNOR2_X1 \myifu/_1693_ ( .A(\myifu/_0764_ ), .B(\myifu/_0306_ ), .ZN(\myifu/_0765_ ) );
XNOR2_X1 \myifu/_1694_ ( .A(\myifu/_0763_ ), .B(\myifu/_0765_ ), .ZN(\myifu/_0766_ ) );
AND3_X1 \myifu/_1695_ ( .A1(\myifu/_0876_ ), .A2(\myifu/_0943_ ), .A3(\myifu/_0929_ ), .ZN(\myifu/_0767_ ) );
OAI22_X1 \myifu/_1696_ ( .A1(\myifu/_0766_ ), .A2(\myifu/_0548_ ), .B1(\myifu/_0567_ ), .B2(\myifu/_0767_ ), .ZN(\myifu/_0768_ ) );
OAI21_X1 \myifu/_1697_ ( .A(\myifu/_0052_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0769_ ) );
AOI21_X1 \myifu/_1698_ ( .A(fanout_net_18 ), .B1(\myifu/_0768_ ), .B2(\myifu/_0769_ ), .ZN(\myifu/_0093_ ) );
AND2_X2 \myifu/_1699_ ( .A1(\myifu/_0757_ ), .A2(\myifu/_0765_ ), .ZN(\myifu/_0770_ ) );
AND3_X2 \myifu/_1700_ ( .A1(\myifu/_0770_ ), .A2(\myifu/_0727_ ), .A3(\myifu/_0745_ ), .ZN(\myifu/_0771_ ) );
AND4_X4 \myifu/_1701_ ( .A1(\myifu/_0656_ ), .A2(\myifu/_0678_ ), .A3(\myifu/_0679_ ), .A4(\myifu/_0730_ ), .ZN(\myifu/_0772_ ) );
OR4_X4 \myifu/_1702_ ( .A1(\myifu/_0718_ ), .A2(\myifu/_0732_ ), .A3(\myifu/_0733_ ), .A4(\myifu/_0736_ ), .ZN(\myifu/_0773_ ) );
OAI21_X2 \myifu/_1703_ ( .A(\myifu/_0771_ ), .B1(\myifu/_0772_ ), .B2(\myifu/_0773_ ), .ZN(\myifu/_0774_ ) );
INV_X1 \myifu/_1704_ ( .A(\myifu/_0754_ ), .ZN(\myifu/_0775_ ) );
OAI21_X1 \myifu/_1705_ ( .A(\myifu/_0775_ ), .B1(\myifu/_0746_ ), .B2(\myifu/_0748_ ), .ZN(\myifu/_0776_ ) );
AND2_X1 \myifu/_1706_ ( .A1(\myifu/_0770_ ), .A2(\myifu/_0776_ ), .ZN(\myifu/_0777_ ) );
NOR3_X1 \myifu/_1707_ ( .A1(\myifu/_0600_ ), .A2(\myifu/_0306_ ), .A3(\myifu/_0039_ ), .ZN(\myifu/_0778_ ) );
AND3_X1 \myifu/_1708_ ( .A1(\myifu/_0765_ ), .A2(\myifu/_0051_ ), .A3(\myifu/_0756_ ), .ZN(\myifu/_0779_ ) );
NOR3_X4 \myifu/_1709_ ( .A1(\myifu/_0777_ ), .A2(\myifu/_0778_ ), .A3(\myifu/_0779_ ), .ZN(\myifu/_0780_ ) );
AND2_X4 \myifu/_1710_ ( .A1(\myifu/_0774_ ), .A2(\myifu/_0780_ ), .ZN(\myifu/_0781_ ) );
BUF_X4 \myifu/_1711_ ( .A(\myifu/_0764_ ), .Z(\myifu/_0782_ ) );
INV_X1 \myifu/_1712_ ( .A(\myifu/_0053_ ), .ZN(\myifu/_0783_ ) );
XNOR2_X1 \myifu/_1713_ ( .A(\myifu/_0782_ ), .B(\myifu/_0783_ ), .ZN(\myifu/_0784_ ) );
INV_X1 \myifu/_1714_ ( .A(\myifu/_0784_ ), .ZN(\myifu/_0785_ ) );
NOR2_X1 \myifu/_1715_ ( .A1(\myifu/_0781_ ), .A2(\myifu/_0785_ ), .ZN(\myifu/_0786_ ) );
AND3_X1 \myifu/_1716_ ( .A1(\myifu/_0774_ ), .A2(\myifu/_0780_ ), .A3(\myifu/_0785_ ), .ZN(\myifu/_0787_ ) );
OR4_X1 \myifu/_1717_ ( .A1(\myifu/_0548_ ), .A2(\myifu/_0786_ ), .A3(\myifu/_0525_ ), .A4(\myifu/_0787_ ), .ZN(\myifu/_0788_ ) );
AOI22_X1 \myifu/_1718_ ( .A1(\myifu/_0531_ ), .A2(\myifu/_0877_ ), .B1(\myifu/_0053_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0789_ ) );
AOI21_X1 \myifu/_1719_ ( .A(fanout_net_18 ), .B1(\myifu/_0788_ ), .B2(\myifu/_0789_ ), .ZN(\myifu/_0094_ ) );
NOR3_X1 \myifu/_1720_ ( .A1(\myifu/_0600_ ), .A2(\myifu/_0783_ ), .A3(\myifu/_0039_ ), .ZN(\myifu/_0790_ ) );
OR2_X1 \myifu/_1721_ ( .A1(\myifu/_0786_ ), .A2(\myifu/_0790_ ), .ZN(\myifu/_0791_ ) );
XNOR2_X1 \myifu/_1722_ ( .A(\myifu/_0782_ ), .B(\myifu/_0041_ ), .ZN(\myifu/_0792_ ) );
INV_X1 \myifu/_1723_ ( .A(\myifu/_0792_ ), .ZN(\myifu/_0793_ ) );
AND2_X1 \myifu/_1724_ ( .A1(\myifu/_0791_ ), .A2(\myifu/_0793_ ), .ZN(\myifu/_0794_ ) );
OAI21_X1 \myifu/_1725_ ( .A(\myifu/_0528_ ), .B1(\myifu/_0791_ ), .B2(\myifu/_0793_ ), .ZN(\myifu/_0795_ ) );
OAI221_X1 \myifu/_1726_ ( .A(\myifu/_0547_ ), .B1(\myifu/_0878_ ), .B2(\myifu/_0571_ ), .C1(\myifu/_0794_ ), .C2(\myifu/_0795_ ), .ZN(\myifu/_0796_ ) );
OAI21_X1 \myifu/_1727_ ( .A(\myifu/_0054_ ), .B1(\myifu/_0236_ ), .B2(\myifu/_0345_ ), .ZN(\myifu/_0797_ ) );
AOI21_X1 \myifu/_1728_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0796_ ), .B2(\myifu/_0797_ ), .ZN(\myifu/_0095_ ) );
OR3_X4 \myifu/_1729_ ( .A1(\myifu/_0781_ ), .A2(\myifu/_0785_ ), .A3(\myifu/_0793_ ), .ZN(\myifu/_0798_ ) );
AND3_X1 \myifu/_1730_ ( .A1(\myifu/_0782_ ), .A2(\myifu/_0053_ ), .A3(\myifu/_0041_ ), .ZN(\myifu/_0799_ ) );
AOI21_X1 \myifu/_1731_ ( .A(\myifu/_0799_ ), .B1(\myifu/_0054_ ), .B2(\myifu/_0782_ ), .ZN(\myifu/_0800_ ) );
AND2_X4 \myifu/_1732_ ( .A1(\myifu/_0798_ ), .A2(\myifu/_0800_ ), .ZN(\myifu/_0801_ ) );
XNOR2_X1 \myifu/_1733_ ( .A(\myifu/_0764_ ), .B(\myifu/_0288_ ), .ZN(\myifu/_0802_ ) );
INV_X1 \myifu/_1734_ ( .A(\myifu/_0802_ ), .ZN(\myifu/_0803_ ) );
OR2_X4 \myifu/_1735_ ( .A1(\myifu/_0801_ ), .A2(\myifu/_0803_ ), .ZN(\myifu/_0804_ ) );
NAND3_X1 \myifu/_1736_ ( .A1(\myifu/_0798_ ), .A2(\myifu/_0800_ ), .A3(\myifu/_0803_ ), .ZN(\myifu/_0805_ ) );
NAND3_X1 \myifu/_1737_ ( .A1(\myifu/_0804_ ), .A2(\myifu/_0567_ ), .A3(\myifu/_0805_ ), .ZN(\myifu/_0806_ ) );
AOI22_X1 \myifu/_1738_ ( .A1(\myifu/_0531_ ), .A2(\myifu/_0879_ ), .B1(\myifu/_0055_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0807_ ) );
AOI21_X1 \myifu/_1739_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0806_ ), .B2(\myifu/_0807_ ), .ZN(\myifu/_0096_ ) );
BUF_X4 \myifu/_1740_ ( .A(\myifu/_0782_ ), .Z(\myifu/_0808_ ) );
NAND2_X1 \myifu/_1741_ ( .A1(\myifu/_0808_ ), .A2(\myifu/_0055_ ), .ZN(\myifu/_0809_ ) );
NAND2_X4 \myifu/_1742_ ( .A1(\myifu/_0804_ ), .A2(\myifu/_0809_ ), .ZN(\myifu/_0810_ ) );
XNOR2_X1 \myifu/_1743_ ( .A(\myifu/_0782_ ), .B(\myifu/_0056_ ), .ZN(\myifu/_0811_ ) );
AND2_X2 \myifu/_1744_ ( .A1(\myifu/_0810_ ), .A2(\myifu/_0811_ ), .ZN(\myifu/_0812_ ) );
OAI21_X1 \myifu/_1745_ ( .A(\myifu/_0528_ ), .B1(\myifu/_0810_ ), .B2(\myifu/_0811_ ), .ZN(\myifu/_0813_ ) );
OAI221_X1 \myifu/_1746_ ( .A(\myifu/_0547_ ), .B1(\myifu/_0880_ ), .B2(\myifu/_0571_ ), .C1(\myifu/_0812_ ), .C2(\myifu/_0813_ ), .ZN(\myifu/_0814_ ) );
OAI21_X1 \myifu/_1747_ ( .A(\myifu/_0056_ ), .B1(\myifu/_0235_ ), .B2(\myifu/_0344_ ), .ZN(\myifu/_0815_ ) );
AOI21_X1 \myifu/_1748_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0814_ ), .B2(\myifu/_0815_ ), .ZN(\myifu/_0097_ ) );
NOR3_X1 \myifu/_1749_ ( .A1(\myifu/_0793_ ), .A2(\myifu/_0803_ ), .A3(\myifu/_0811_ ), .ZN(\myifu/_0816_ ) );
NAND3_X1 \myifu/_1750_ ( .A1(\myifu/_0771_ ), .A2(\myifu/_0784_ ), .A3(\myifu/_0816_ ), .ZN(\myifu/_0817_ ) );
AOI21_X4 \myifu/_1751_ ( .A(\myifu/_0817_ ), .B1(\myifu/_0731_ ), .B2(\myifu/_0737_ ), .ZN(\myifu/_0818_ ) );
OR3_X1 \myifu/_1752_ ( .A1(\myifu/_0800_ ), .A2(\myifu/_0803_ ), .A3(\myifu/_0811_ ), .ZN(\myifu/_0819_ ) );
OAI21_X1 \myifu/_1753_ ( .A(\myifu/_0782_ ), .B1(\myifu/_0055_ ), .B2(\myifu/_0056_ ), .ZN(\myifu/_0820_ ) );
NAND2_X1 \myifu/_1754_ ( .A1(\myifu/_0816_ ), .A2(\myifu/_0784_ ), .ZN(\myifu/_0821_ ) );
OAI211_X2 \myifu/_1755_ ( .A(\myifu/_0819_ ), .B(\myifu/_0820_ ), .C1(\myifu/_0780_ ), .C2(\myifu/_0821_ ), .ZN(\myifu/_0822_ ) );
XOR2_X1 \myifu/_1756_ ( .A(\myifu/_0782_ ), .B(\myifu/_0057_ ), .Z(\myifu/_0823_ ) );
OR3_X1 \myifu/_1757_ ( .A1(\myifu/_0818_ ), .A2(\myifu/_0822_ ), .A3(\myifu/_0823_ ), .ZN(\myifu/_0824_ ) );
OAI21_X1 \myifu/_1758_ ( .A(\myifu/_0823_ ), .B1(\myifu/_0818_ ), .B2(\myifu/_0822_ ), .ZN(\myifu/_0825_ ) );
NAND3_X1 \myifu/_1759_ ( .A1(\myifu/_0824_ ), .A2(\myifu/_0567_ ), .A3(\myifu/_0825_ ), .ZN(\myifu/_0826_ ) );
AOI22_X1 \myifu/_1760_ ( .A1(\myifu/_0531_ ), .A2(\myifu/_0881_ ), .B1(\myifu/_0057_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0827_ ) );
AOI21_X1 \myifu/_1761_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0826_ ), .B2(\myifu/_0827_ ), .ZN(\myifu/_0098_ ) );
NAND2_X1 \myifu/_1762_ ( .A1(\myifu/_0808_ ), .A2(\myifu/_0057_ ), .ZN(\myifu/_0828_ ) );
AND2_X1 \myifu/_1763_ ( .A1(\myifu/_0825_ ), .A2(\myifu/_0828_ ), .ZN(\myifu/_0829_ ) );
XNOR2_X1 \myifu/_1764_ ( .A(\myifu/_0782_ ), .B(\myifu/_0285_ ), .ZN(\myifu/_0830_ ) );
XNOR2_X1 \myifu/_1765_ ( .A(\myifu/_0829_ ), .B(\myifu/_0830_ ), .ZN(\myifu/_0831_ ) );
AND3_X1 \myifu/_1766_ ( .A1(\myifu/_0882_ ), .A2(\myifu/_0943_ ), .A3(\myifu/_0929_ ), .ZN(\myifu/_0832_ ) );
OAI22_X1 \myifu/_1767_ ( .A1(\myifu/_0831_ ), .A2(\myifu/_0548_ ), .B1(\myifu/_0567_ ), .B2(\myifu/_0832_ ), .ZN(\myifu/_0833_ ) );
OAI21_X1 \myifu/_1768_ ( .A(\myifu/_0058_ ), .B1(\myifu/_0235_ ), .B2(\myifu/_0344_ ), .ZN(\myifu/_0834_ ) );
AOI21_X1 \myifu/_1769_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0833_ ), .B2(\myifu/_0834_ ), .ZN(\myifu/_0099_ ) );
NOR2_X1 \myifu/_1770_ ( .A1(\myifu/_0818_ ), .A2(\myifu/_0822_ ), .ZN(\myifu/_0835_ ) );
INV_X1 \myifu/_1771_ ( .A(\myifu/_0835_ ), .ZN(\myifu/_0836_ ) );
AND2_X1 \myifu/_1772_ ( .A1(\myifu/_0823_ ), .A2(\myifu/_0830_ ), .ZN(\myifu/_0837_ ) );
AND2_X4 \myifu/_1773_ ( .A1(\myifu/_0836_ ), .A2(\myifu/_0837_ ), .ZN(\myifu/_0838_ ) );
OAI21_X1 \myifu/_1774_ ( .A(\myifu/_0808_ ), .B1(\myifu/_0057_ ), .B2(\myifu/_0058_ ), .ZN(\myifu/_0839_ ) );
INV_X1 \myifu/_1775_ ( .A(\myifu/_0839_ ), .ZN(\myifu/_0840_ ) );
INV_X1 \myifu/_1776_ ( .A(\myifu/_0059_ ), .ZN(\myifu/_0841_ ) );
XNOR2_X1 \myifu/_1777_ ( .A(\myifu/_0808_ ), .B(\myifu/_0841_ ), .ZN(\myifu/_0842_ ) );
OR3_X1 \myifu/_1778_ ( .A1(\myifu/_0838_ ), .A2(\myifu/_0840_ ), .A3(\myifu/_0842_ ), .ZN(\myifu/_0843_ ) );
OAI21_X4 \myifu/_1779_ ( .A(\myifu/_0842_ ), .B1(\myifu/_0838_ ), .B2(\myifu/_0840_ ), .ZN(\myifu/_0844_ ) );
NAND3_X1 \myifu/_1780_ ( .A1(\myifu/_0843_ ), .A2(\myifu/_0567_ ), .A3(\myifu/_0844_ ), .ZN(\myifu/_0845_ ) );
AOI22_X1 \myifu/_1781_ ( .A1(\myifu/_0531_ ), .A2(\myifu/_0883_ ), .B1(\myifu/_0059_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0846_ ) );
AOI21_X1 \myifu/_1782_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0845_ ), .B2(\myifu/_0846_ ), .ZN(\myifu/_0100_ ) );
AND2_X1 \myifu/_1783_ ( .A1(\myifu/_0808_ ), .A2(\myifu/_0059_ ), .ZN(\myifu/_0847_ ) );
INV_X1 \myifu/_1784_ ( .A(\myifu/_0847_ ), .ZN(\myifu/_0848_ ) );
AND2_X4 \myifu/_1785_ ( .A1(\myifu/_0844_ ), .A2(\myifu/_0848_ ), .ZN(\myifu/_0849_ ) );
XNOR2_X1 \myifu/_1786_ ( .A(\myifu/_0782_ ), .B(\myifu/_0333_ ), .ZN(\myifu/_0850_ ) );
XNOR2_X2 \myifu/_1787_ ( .A(\myifu/_0849_ ), .B(\myifu/_0850_ ), .ZN(\myifu/_0851_ ) );
MUX2_X2 \myifu/_1788_ ( .A(\myifu/_0884_ ), .B(\myifu/_0851_ ), .S(\myifu/_0528_ ), .Z(\myifu/_0852_ ) );
NAND2_X2 \myifu/_1789_ ( .A1(\myifu/_0852_ ), .A2(\myifu/_0547_ ), .ZN(\myifu/_0853_ ) );
OAI211_X2 \myifu/_1790_ ( .A(\myifu/_0853_ ), .B(\myifu/_0343_ ), .C1(\myifu/_0333_ ), .C2(\myifu/_0547_ ), .ZN(\myifu/_0101_ ) );
AND2_X1 \myifu/_1791_ ( .A1(\myifu/_0842_ ), .A2(\myifu/_0850_ ), .ZN(\myifu/_0854_ ) );
OAI211_X2 \myifu/_1792_ ( .A(\myifu/_0837_ ), .B(\myifu/_0854_ ), .C1(\myifu/_0818_ ), .C2(\myifu/_0822_ ), .ZN(\myifu/_0855_ ) );
AOI221_X4 \myifu/_1793_ ( .A(\myifu/_0039_ ), .B1(\myifu/_0841_ ), .B2(\myifu/_0333_ ), .C1(\myifu/_0562_ ), .C2(\myifu/_0587_ ), .ZN(\myifu/_0856_ ) );
AOI21_X1 \myifu/_1794_ ( .A(\myifu/_0856_ ), .B1(\myifu/_0854_ ), .B2(\myifu/_0840_ ), .ZN(\myifu/_0857_ ) );
NAND2_X2 \myifu/_1795_ ( .A1(\myifu/_0855_ ), .A2(\myifu/_0857_ ), .ZN(\myifu/_0205_ ) );
XNOR2_X1 \myifu/_1796_ ( .A(\myifu/_0808_ ), .B(\myifu/_0328_ ), .ZN(\myifu/_0206_ ) );
AOI211_X4 \myifu/_1797_ ( .A(\myifu/_0548_ ), .B(\myifu/_0524_ ), .C1(\myifu/_0205_ ), .C2(\myifu/_0206_ ), .ZN(\myifu/_0207_ ) );
OAI21_X1 \myifu/_1798_ ( .A(\myifu/_0207_ ), .B1(\myifu/_0205_ ), .B2(\myifu/_0206_ ), .ZN(\myifu/_0208_ ) );
AOI221_X4 \myifu/_1799_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0061_ ), .B2(\myifu/_0524_ ), .C1(\myifu/_0531_ ), .C2(\myifu/_0885_ ), .ZN(\myifu/_0209_ ) );
NAND2_X1 \myifu/_1800_ ( .A1(\myifu/_0208_ ), .A2(\myifu/_0209_ ), .ZN(\myifu/_0102_ ) );
NAND2_X1 \myifu/_1801_ ( .A1(\myifu/_0205_ ), .A2(\myifu/_0206_ ), .ZN(\myifu/_0210_ ) );
NAND2_X1 \myifu/_1802_ ( .A1(\myifu/_0808_ ), .A2(\myifu/_0061_ ), .ZN(\myifu/_0211_ ) );
AND2_X1 \myifu/_1803_ ( .A1(\myifu/_0210_ ), .A2(\myifu/_0211_ ), .ZN(\myifu/_0212_ ) );
XNOR2_X1 \myifu/_1804_ ( .A(\myifu/_0808_ ), .B(\myifu/_0334_ ), .ZN(\myifu/_0213_ ) );
AOI21_X1 \myifu/_1805_ ( .A(\myifu/_0548_ ), .B1(\myifu/_0212_ ), .B2(\myifu/_0213_ ), .ZN(\myifu/_0214_ ) );
OAI21_X1 \myifu/_1806_ ( .A(\myifu/_0214_ ), .B1(\myifu/_0212_ ), .B2(\myifu/_0213_ ), .ZN(\myifu/_0215_ ) );
OAI211_X2 \myifu/_1807_ ( .A(\myifu/_0215_ ), .B(\myifu/_0547_ ), .C1(\myifu/_0887_ ), .C2(\myifu/_0571_ ), .ZN(\myifu/_0216_ ) );
OAI21_X1 \myifu/_1808_ ( .A(\myifu/_0062_ ), .B1(\myifu/_0235_ ), .B2(\myifu/_0344_ ), .ZN(\myifu/_0217_ ) );
AOI21_X1 \myifu/_1809_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0216_ ), .B2(\myifu/_0217_ ), .ZN(\myifu/_0103_ ) );
NAND3_X2 \myifu/_1810_ ( .A1(\myifu/_0205_ ), .A2(\myifu/_0206_ ), .A3(\myifu/_0213_ ), .ZN(\myifu/_0218_ ) );
OAI21_X1 \myifu/_1811_ ( .A(\myifu/_0808_ ), .B1(\myifu/_0061_ ), .B2(\myifu/_0062_ ), .ZN(\myifu/_0219_ ) );
XNOR2_X1 \myifu/_1812_ ( .A(\myifu/_0808_ ), .B(\myifu/_0063_ ), .ZN(\myifu/_0220_ ) );
AND3_X1 \myifu/_1813_ ( .A1(\myifu/_0218_ ), .A2(\myifu/_0219_ ), .A3(\myifu/_0220_ ), .ZN(\myifu/_0221_ ) );
AOI21_X1 \myifu/_1814_ ( .A(\myifu/_0220_ ), .B1(\myifu/_0218_ ), .B2(\myifu/_0219_ ), .ZN(\myifu/_0222_ ) );
OR4_X2 \myifu/_1815_ ( .A1(\myifu/_0548_ ), .A2(\myifu/_0221_ ), .A3(\myifu/_0222_ ), .A4(\myifu/_0524_ ), .ZN(\myifu/_0223_ ) );
AOI22_X1 \myifu/_1816_ ( .A1(\myifu/_0531_ ), .A2(\myifu/_0888_ ), .B1(\myifu/_0063_ ), .B2(\myifu/_0525_ ), .ZN(\myifu/_0224_ ) );
AOI21_X1 \myifu/_1817_ ( .A(\myifu/_0930_ ), .B1(\myifu/_0223_ ), .B2(\myifu/_0224_ ), .ZN(\myifu/_0104_ ) );
AND2_X1 \myifu/_1818_ ( .A1(\myifu/_0351_ ), .A2(\myifu/_0944_ ), .ZN(\myifu/_0225_ ) );
INV_X1 \myifu/_1819_ ( .A(\myifu/_0225_ ), .ZN(\myifu/_0226_ ) );
NOR2_X1 \myifu/_1820_ ( .A1(\myifu/_0935_ ), .A2(\myifu/_0972_ ), .ZN(\myifu/_0227_ ) );
NOR2_X1 \myifu/_1821_ ( .A1(\myifu/_0226_ ), .A2(\myifu/_0227_ ), .ZN(\myifu/_0228_ ) );
AOI211_X4 \myifu/_1822_ ( .A(\myifu/_0930_ ), .B(\myifu/_0228_ ), .C1(\myifu/_0373_ ), .C2(\myifu/_0226_ ), .ZN(\myifu/_0105_ ) );
AOI21_X1 \myifu/_1823_ ( .A(\myifu/_0365_ ), .B1(\myifu/_0355_ ), .B2(\myifu/_0071_ ), .ZN(\myifu/_0229_ ) );
OAI21_X1 \myifu/_1824_ ( .A(\myifu/_0369_ ), .B1(\myifu/_0357_ ), .B2(\myifu/_0358_ ), .ZN(\myifu/_0230_ ) );
NOR2_X1 \myifu/_1825_ ( .A1(\myifu/_0229_ ), .A2(\myifu/_0230_ ), .ZN(\myifu/_0231_ ) );
OAI21_X1 \myifu/_1826_ ( .A(\myifu/_0343_ ), .B1(\myifu/_0231_ ), .B2(\myifu/_0974_ ), .ZN(\myifu/_0232_ ) );
NOR3_X1 \myifu/_1827_ ( .A1(\myifu/_0229_ ), .A2(\myifu/_0024_ ), .A3(\myifu/_0230_ ), .ZN(\myifu/_0233_ ) );
NOR2_X1 \myifu/_1828_ ( .A1(\myifu/_0232_ ), .A2(\myifu/_0233_ ), .ZN(\myifu/_0138_ ) );
DFF_X1 \myifu/_1829_ ( .D(\myifu/_1031_ ), .CK(clock ), .Q(\IF_ID_pc [0] ), .QN(\myifu/_0005_ ) );
DFF_X1 \myifu/_1830_ ( .D(\myifu/_0000_ ), .CK(clock ), .Q(\myifu/state [0] ), .QN(\myifu/_1027_ ) );
DFF_X1 \myifu/_1831_ ( .D(\myifu/_0001_ ), .CK(clock ), .Q(\myifu/state [1] ), .QN(\myifu/_1028_ ) );
DFF_X1 \myifu/_1832_ ( .D(\myifu/_0002_ ), .CK(clock ), .Q(\myifu/state [2] ), .QN(\myifu/_0003_ ) );
DFF_X1 \myifu/_1833_ ( .D(\myifu/_1032_ ), .CK(clock ), .Q(\IF_ID_pc [1] ), .QN(\myifu/_0006_ ) );
DFF_X1 \myifu/_1834_ ( .D(\myifu/_1033_ ), .CK(clock ), .Q(\IF_ID_pc [2] ), .QN(\myifu/_1026_ ) );
DFF_X1 \myifu/_1835_ ( .D(\myifu/_1034_ ), .CK(clock ), .Q(\araddr_IFU [3] ), .QN(\myifu/_1025_ ) );
DFF_X1 \myifu/_1836_ ( .D(\myifu/_1035_ ), .CK(clock ), .Q(\araddr_IFU [4] ), .QN(\myifu/_1024_ ) );
DFF_X1 \myifu/_1837_ ( .D(\myifu/_1036_ ), .CK(clock ), .Q(\araddr_IFU [5] ), .QN(\myifu/_1023_ ) );
DFF_X1 \myifu/_1838_ ( .D(\myifu/_1037_ ), .CK(clock ), .Q(\araddr_IFU [6] ), .QN(\myifu/_1022_ ) );
DFF_X1 \myifu/_1839_ ( .D(\myifu/_1038_ ), .CK(clock ), .Q(\araddr_IFU [7] ), .QN(\myifu/_1021_ ) );
DFF_X1 \myifu/_1840_ ( .D(\myifu/_1039_ ), .CK(clock ), .Q(\araddr_IFU [8] ), .QN(\myifu/_1020_ ) );
DFF_X1 \myifu/_1841_ ( .D(\myifu/_1040_ ), .CK(clock ), .Q(\araddr_IFU [9] ), .QN(\myifu/_1019_ ) );
DFF_X1 \myifu/_1842_ ( .D(\myifu/_1041_ ), .CK(clock ), .Q(\araddr_IFU [10] ), .QN(\myifu/_1018_ ) );
DFF_X1 \myifu/_1843_ ( .D(\myifu/_1042_ ), .CK(clock ), .Q(\araddr_IFU [11] ), .QN(\myifu/_1017_ ) );
DFF_X1 \myifu/_1844_ ( .D(\myifu/_1043_ ), .CK(clock ), .Q(\araddr_IFU [12] ), .QN(\myifu/_1016_ ) );
DFF_X1 \myifu/_1845_ ( .D(\myifu/_1044_ ), .CK(clock ), .Q(\araddr_IFU [13] ), .QN(\myifu/_1015_ ) );
DFF_X1 \myifu/_1846_ ( .D(\myifu/_1045_ ), .CK(clock ), .Q(\araddr_IFU [14] ), .QN(\myifu/_1014_ ) );
DFF_X1 \myifu/_1847_ ( .D(\myifu/_1046_ ), .CK(clock ), .Q(\araddr_IFU [15] ), .QN(\myifu/_1013_ ) );
DFF_X1 \myifu/_1848_ ( .D(\myifu/_1047_ ), .CK(clock ), .Q(\araddr_IFU [16] ), .QN(\myifu/_1012_ ) );
DFF_X1 \myifu/_1849_ ( .D(\myifu/_1048_ ), .CK(clock ), .Q(\araddr_IFU [17] ), .QN(\myifu/_1011_ ) );
DFF_X1 \myifu/_1850_ ( .D(\myifu/_1049_ ), .CK(clock ), .Q(\araddr_IFU [18] ), .QN(\myifu/_0019_ ) );
DFF_X1 \myifu/_1851_ ( .D(\myifu/_1050_ ), .CK(clock ), .Q(\araddr_IFU [19] ), .QN(\myifu/_1010_ ) );
DFF_X1 \myifu/_1852_ ( .D(\myifu/_1051_ ), .CK(clock ), .Q(\araddr_IFU [20] ), .QN(\myifu/_1009_ ) );
DFF_X1 \myifu/_1853_ ( .D(\myifu/_1052_ ), .CK(clock ), .Q(\araddr_IFU [21] ), .QN(\myifu/_1008_ ) );
DFF_X1 \myifu/_1854_ ( .D(\myifu/_1053_ ), .CK(clock ), .Q(\araddr_IFU [22] ), .QN(\myifu/_0020_ ) );
DFF_X1 \myifu/_1855_ ( .D(\myifu/_1054_ ), .CK(clock ), .Q(\araddr_IFU [23] ), .QN(\myifu/_1007_ ) );
DFF_X1 \myifu/_1856_ ( .D(\myifu/_1055_ ), .CK(clock ), .Q(\araddr_IFU [24] ), .QN(\myifu/_1006_ ) );
DFF_X1 \myifu/_1857_ ( .D(\myifu/_1056_ ), .CK(clock ), .Q(\araddr_IFU [25] ), .QN(\myifu/_1005_ ) );
DFF_X1 \myifu/_1858_ ( .D(\myifu/_1057_ ), .CK(clock ), .Q(\araddr_IFU [26] ), .QN(\myifu/_1004_ ) );
DFF_X1 \myifu/_1859_ ( .D(\myifu/_1058_ ), .CK(clock ), .Q(\araddr_IFU [27] ), .QN(\myifu/_1003_ ) );
DFF_X1 \myifu/_1860_ ( .D(\myifu/_1059_ ), .CK(clock ), .Q(\araddr_IFU [28] ), .QN(\myifu/_1002_ ) );
DFF_X1 \myifu/_1861_ ( .D(\myifu/_1060_ ), .CK(clock ), .Q(\araddr_IFU [29] ), .QN(\myifu/_1001_ ) );
DFF_X1 \myifu/_1862_ ( .D(\myifu/_1061_ ), .CK(clock ), .Q(\araddr_IFU [30] ), .QN(\myifu/_1000_ ) );
DFF_X1 \myifu/_1863_ ( .D(\myifu/_1062_ ), .CK(clock ), .Q(\araddr_IFU [31] ), .QN(\myifu/_0999_ ) );
DFF_X1 \myifu/_1864_ ( .D(\myifu/_1063_ ), .CK(clock ), .Q(\myifu/tmp_offset [2] ), .QN(\myifu/_0998_ ) );
DFF_X1 \myifu/_1865_ ( .D(\myifu/_1064_ ), .CK(clock ), .Q(\IF_ID_inst [0] ), .QN(\myifu/_0997_ ) );
DFF_X1 \myifu/_1866_ ( .D(\myifu/_1065_ ), .CK(clock ), .Q(\IF_ID_inst [1] ), .QN(\myifu/_0996_ ) );
DFF_X1 \myifu/_1867_ ( .D(\myifu/_1066_ ), .CK(clock ), .Q(\IF_ID_inst [2] ), .QN(\myifu/_0995_ ) );
DFF_X1 \myifu/_1868_ ( .D(\myifu/_1067_ ), .CK(clock ), .Q(\IF_ID_inst [3] ), .QN(\myifu/_0994_ ) );
DFF_X1 \myifu/_1869_ ( .D(\myifu/_1068_ ), .CK(clock ), .Q(\IF_ID_inst [4] ), .QN(\myifu/_0993_ ) );
DFF_X1 \myifu/_1870_ ( .D(\myifu/_1069_ ), .CK(clock ), .Q(\IF_ID_inst [5] ), .QN(\myifu/_0992_ ) );
DFF_X1 \myifu/_1871_ ( .D(\myifu/_1070_ ), .CK(clock ), .Q(\IF_ID_inst [6] ), .QN(\myifu/_0991_ ) );
DFF_X1 \myifu/_1872_ ( .D(\myifu/_1071_ ), .CK(clock ), .Q(\IF_ID_inst [7] ), .QN(\myifu/_0017_ ) );
DFF_X1 \myifu/_1873_ ( .D(\myifu/_1072_ ), .CK(clock ), .Q(\IF_ID_inst [8] ), .QN(\myifu/_0007_ ) );
DFF_X1 \myifu/_1874_ ( .D(\myifu/_1073_ ), .CK(clock ), .Q(\IF_ID_inst [9] ), .QN(\myifu/_0008_ ) );
DFF_X1 \myifu/_1875_ ( .D(\myifu/_1074_ ), .CK(clock ), .Q(\IF_ID_inst [10] ), .QN(\myifu/_0009_ ) );
DFF_X1 \myifu/_1876_ ( .D(\myifu/_1075_ ), .CK(clock ), .Q(\IF_ID_inst [11] ), .QN(\myifu/_0010_ ) );
DFF_X1 \myifu/_1877_ ( .D(\myifu/_1076_ ), .CK(clock ), .Q(\IF_ID_inst [12] ), .QN(\myifu/_0990_ ) );
DFF_X1 \myifu/_1878_ ( .D(\myifu/_1077_ ), .CK(clock ), .Q(\IF_ID_inst [13] ), .QN(\myifu/_0989_ ) );
DFF_X1 \myifu/_1879_ ( .D(\myifu/_1078_ ), .CK(clock ), .Q(\IF_ID_inst [14] ), .QN(\myifu/_0988_ ) );
DFF_X1 \myifu/_1880_ ( .D(\myifu/_1079_ ), .CK(clock ), .Q(\IF_ID_inst [15] ), .QN(\myifu/_0987_ ) );
DFF_X1 \myifu/_1881_ ( .D(\myifu/_1080_ ), .CK(clock ), .Q(\IF_ID_inst [16] ), .QN(\myifu/_0986_ ) );
DFF_X1 \myifu/_1882_ ( .D(\myifu/_1081_ ), .CK(clock ), .Q(\IF_ID_inst [17] ), .QN(\myifu/_0985_ ) );
DFF_X1 \myifu/_1883_ ( .D(\myifu/_1082_ ), .CK(clock ), .Q(\IF_ID_inst [18] ), .QN(\myifu/_0984_ ) );
DFF_X1 \myifu/_1884_ ( .D(\myifu/_1083_ ), .CK(clock ), .Q(\IF_ID_inst [19] ), .QN(\myifu/_0983_ ) );
DFF_X1 \myifu/_1885_ ( .D(\myifu/_1084_ ), .CK(clock ), .Q(\IF_ID_inst [20] ), .QN(\myifu/_0982_ ) );
DFF_X1 \myifu/_1886_ ( .D(\myifu/_1085_ ), .CK(clock ), .Q(\IF_ID_inst [21] ), .QN(\myifu/_0981_ ) );
DFF_X1 \myifu/_1887_ ( .D(\myifu/_1086_ ), .CK(clock ), .Q(\IF_ID_inst [22] ), .QN(\myifu/_0980_ ) );
DFF_X1 \myifu/_1888_ ( .D(\myifu/_1087_ ), .CK(clock ), .Q(\IF_ID_inst [23] ), .QN(\myifu/_0979_ ) );
DFF_X1 \myifu/_1889_ ( .D(\myifu/_1088_ ), .CK(clock ), .Q(\IF_ID_inst [24] ), .QN(\myifu/_0978_ ) );
DFF_X1 \myifu/_1890_ ( .D(\myifu/_1089_ ), .CK(clock ), .Q(\IF_ID_inst [25] ), .QN(\myifu/_0011_ ) );
DFF_X1 \myifu/_1891_ ( .D(\myifu/_1090_ ), .CK(clock ), .Q(\IF_ID_inst [26] ), .QN(\myifu/_0012_ ) );
DFF_X1 \myifu/_1892_ ( .D(\myifu/_1091_ ), .CK(clock ), .Q(\IF_ID_inst [27] ), .QN(\myifu/_0013_ ) );
DFF_X1 \myifu/_1893_ ( .D(\myifu/_1092_ ), .CK(clock ), .Q(\IF_ID_inst [28] ), .QN(\myifu/_0014_ ) );
DFF_X1 \myifu/_1894_ ( .D(\myifu/_1093_ ), .CK(clock ), .Q(\IF_ID_inst [29] ), .QN(\myifu/_0015_ ) );
DFF_X1 \myifu/_1895_ ( .D(\myifu/_1094_ ), .CK(clock ), .Q(\IF_ID_inst [30] ), .QN(\myifu/_0016_ ) );
DFF_X1 \myifu/_1896_ ( .D(\myifu/_1095_ ), .CK(clock ), .Q(\myifu/pred_jump ), .QN(\myifu/_0018_ ) );
DFF_X1 \myifu/_1897_ ( .D(\myifu/_1096_ ), .CK(clock ), .Q(\myifu/valid_in ), .QN(\myifu/_0977_ ) );
DFF_X1 \myifu/_1898_ ( .D(\myifu/_1097_ ), .CK(clock ), .Q(check_assert ), .QN(\myifu/_0976_ ) );
LOGIC1_X1 \myifu/_1899_ ( .Z(\myifu/_1029_ ) );
LOGIC0_X1 \myifu/_1900_ ( .Z(\myifu/_1030_ ) );
BUF_X1 \myifu/_1901_ ( .A(\myifu/_1030_ ), .Z(\araddr_IFU [0] ) );
BUF_X1 \myifu/_1902_ ( .A(\myifu/_1030_ ), .Z(\araddr_IFU [1] ) );
BUF_X1 \myifu/_1903_ ( .A(\myifu/_1030_ ), .Z(\araddr_IFU [2] ) );
BUF_X1 \myifu/_1904_ ( .A(\myifu/_1029_ ), .Z(\arburst_IFU [0] ) );
BUF_X1 \myifu/_1905_ ( .A(\myifu/_1030_ ), .Z(\arburst_IFU [1] ) );
BUF_X1 \myifu/_1906_ ( .A(\myifu/_1029_ ), .Z(\arid_IFU [0] ) );
BUF_X1 \myifu/_1907_ ( .A(\myifu/_1030_ ), .Z(\arid_IFU [1] ) );
BUF_X1 \myifu/_1908_ ( .A(\myifu/_1030_ ), .Z(\arid_IFU [2] ) );
BUF_X1 \myifu/_1909_ ( .A(\myifu/_1030_ ), .Z(\arid_IFU [3] ) );
BUF_X1 \myifu/_1910_ ( .A(\myifu/_1029_ ), .Z(\arlen_IFU [0] ) );
BUF_X1 \myifu/_1911_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [1] ) );
BUF_X1 \myifu/_1912_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [2] ) );
BUF_X1 \myifu/_1913_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [3] ) );
BUF_X1 \myifu/_1914_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [4] ) );
BUF_X1 \myifu/_1915_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [5] ) );
BUF_X1 \myifu/_1916_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [6] ) );
BUF_X1 \myifu/_1917_ ( .A(\myifu/_1030_ ), .Z(\arlen_IFU [7] ) );
BUF_X1 \myifu/_1918_ ( .A(\myifu/_1030_ ), .Z(\arsize_IFU [0] ) );
BUF_X1 \myifu/_1919_ ( .A(\myifu/_1029_ ), .Z(\arsize_IFU [1] ) );
BUF_X1 \myifu/_1920_ ( .A(\myifu/_1030_ ), .Z(\arsize_IFU [2] ) );
BUF_X1 \myifu/_1921_ ( .A(\myifu/pred_jump ), .Z(\IF_ID_inst [31] ) );
BUF_X1 \myifu/_1922_ ( .A(\araddr_IFU [3] ), .Z(\IF_ID_pc [3] ) );
BUF_X1 \myifu/_1923_ ( .A(\araddr_IFU [4] ), .Z(\IF_ID_pc [4] ) );
BUF_X1 \myifu/_1924_ ( .A(\araddr_IFU [5] ), .Z(\IF_ID_pc [5] ) );
BUF_X1 \myifu/_1925_ ( .A(\araddr_IFU [6] ), .Z(\IF_ID_pc [6] ) );
BUF_X1 \myifu/_1926_ ( .A(\araddr_IFU [7] ), .Z(\IF_ID_pc [7] ) );
BUF_X1 \myifu/_1927_ ( .A(\araddr_IFU [8] ), .Z(\IF_ID_pc [8] ) );
BUF_X1 \myifu/_1928_ ( .A(\araddr_IFU [9] ), .Z(\IF_ID_pc [9] ) );
BUF_X1 \myifu/_1929_ ( .A(\araddr_IFU [10] ), .Z(\IF_ID_pc [10] ) );
BUF_X1 \myifu/_1930_ ( .A(\araddr_IFU [11] ), .Z(\IF_ID_pc [11] ) );
BUF_X1 \myifu/_1931_ ( .A(\araddr_IFU [12] ), .Z(\IF_ID_pc [12] ) );
BUF_X1 \myifu/_1932_ ( .A(\araddr_IFU [13] ), .Z(\IF_ID_pc [13] ) );
BUF_X1 \myifu/_1933_ ( .A(\araddr_IFU [14] ), .Z(\IF_ID_pc [14] ) );
BUF_X1 \myifu/_1934_ ( .A(\araddr_IFU [15] ), .Z(\IF_ID_pc [15] ) );
BUF_X1 \myifu/_1935_ ( .A(\araddr_IFU [16] ), .Z(\IF_ID_pc [16] ) );
BUF_X1 \myifu/_1936_ ( .A(\araddr_IFU [17] ), .Z(\IF_ID_pc [17] ) );
BUF_X1 \myifu/_1937_ ( .A(\araddr_IFU [18] ), .Z(\IF_ID_pc [18] ) );
BUF_X1 \myifu/_1938_ ( .A(\araddr_IFU [19] ), .Z(\IF_ID_pc [19] ) );
BUF_X1 \myifu/_1939_ ( .A(\araddr_IFU [20] ), .Z(\IF_ID_pc [20] ) );
BUF_X1 \myifu/_1940_ ( .A(\araddr_IFU [21] ), .Z(\IF_ID_pc [21] ) );
BUF_X1 \myifu/_1941_ ( .A(\araddr_IFU [22] ), .Z(\IF_ID_pc [22] ) );
BUF_X1 \myifu/_1942_ ( .A(\araddr_IFU [23] ), .Z(\IF_ID_pc [23] ) );
BUF_X1 \myifu/_1943_ ( .A(\araddr_IFU [24] ), .Z(\IF_ID_pc [24] ) );
BUF_X1 \myifu/_1944_ ( .A(\araddr_IFU [25] ), .Z(\IF_ID_pc [25] ) );
BUF_X1 \myifu/_1945_ ( .A(\araddr_IFU [26] ), .Z(\IF_ID_pc [26] ) );
BUF_X1 \myifu/_1946_ ( .A(\araddr_IFU [27] ), .Z(\IF_ID_pc [27] ) );
BUF_X1 \myifu/_1947_ ( .A(\araddr_IFU [28] ), .Z(\IF_ID_pc [28] ) );
BUF_X1 \myifu/_1948_ ( .A(\araddr_IFU [29] ), .Z(\IF_ID_pc [29] ) );
BUF_X1 \myifu/_1949_ ( .A(\araddr_IFU [30] ), .Z(\IF_ID_pc [30] ) );
BUF_X1 \myifu/_1950_ ( .A(\araddr_IFU [31] ), .Z(\IF_ID_pc [31] ) );
BUF_X1 \myifu/_1951_ ( .A(\myifu/_1030_ ), .Z(\myifu/tmp_offset [0] ) );
BUF_X1 \myifu/_1952_ ( .A(\myifu/_1030_ ), .Z(\myifu/tmp_offset [1] ) );
BUF_X1 \myifu/_1953_ ( .A(reset ), .Z(\myifu/_0930_ ) );
BUF_X1 \myifu/_1954_ ( .A(stall_quest_fencei ), .Z(\myifu/_0941_ ) );
BUF_X1 \myifu/_1955_ ( .A(\myifu/state [0] ), .Z(\myifu/_0942_ ) );
BUF_X1 \myifu/_1956_ ( .A(\myifu/_0072_ ), .Z(arvalid_IFU ) );
BUF_X1 \myifu/_1957_ ( .A(\pc_jump [0] ), .Z(\myifu/_0864_ ) );
BUF_X1 \myifu/_1958_ ( .A(\IF_ID_pc [0] ), .Z(\myifu/_0861_ ) );
BUF_X1 \myifu/_1959_ ( .A(\pc_jump [1] ), .Z(\myifu/_0875_ ) );
BUF_X1 \myifu/_1960_ ( .A(\IF_ID_pc [1] ), .Z(\myifu/_0862_ ) );
BUF_X1 \myifu/_1961_ ( .A(\pc_jump [2] ), .Z(\myifu/_0886_ ) );
BUF_X1 \myifu/_1962_ ( .A(\IF_ID_pc [2] ), .Z(\myifu/_0863_ ) );
BUF_X1 \myifu/_1963_ ( .A(\pc_jump [3] ), .Z(\myifu/_0889_ ) );
BUF_X1 \myifu/_1964_ ( .A(\araddr_IFU [3] ), .Z(\myifu/_0064_ ) );
BUF_X1 \myifu/_1965_ ( .A(\pc_jump [4] ), .Z(\myifu/_0890_ ) );
BUF_X1 \myifu/_1966_ ( .A(\araddr_IFU [4] ), .Z(\myifu/_0065_ ) );
BUF_X1 \myifu/_1967_ ( .A(\pc_jump [5] ), .Z(\myifu/_0891_ ) );
BUF_X1 \myifu/_1968_ ( .A(\araddr_IFU [5] ), .Z(\myifu/_0066_ ) );
BUF_X1 \myifu/_1969_ ( .A(\pc_jump [6] ), .Z(\myifu/_0892_ ) );
BUF_X1 \myifu/_1970_ ( .A(\araddr_IFU [6] ), .Z(\myifu/_0067_ ) );
BUF_X1 \myifu/_1971_ ( .A(\pc_jump [7] ), .Z(\myifu/_0893_ ) );
BUF_X1 \myifu/_1972_ ( .A(\araddr_IFU [7] ), .Z(\myifu/_0068_ ) );
BUF_X1 \myifu/_1973_ ( .A(\pc_jump [8] ), .Z(\myifu/_0894_ ) );
BUF_X1 \myifu/_1974_ ( .A(\araddr_IFU [8] ), .Z(\myifu/_0069_ ) );
BUF_X1 \myifu/_1975_ ( .A(\pc_jump [9] ), .Z(\myifu/_0895_ ) );
BUF_X1 \myifu/_1976_ ( .A(\araddr_IFU [9] ), .Z(\myifu/_0070_ ) );
BUF_X1 \myifu/_1977_ ( .A(\pc_jump [10] ), .Z(\myifu/_0865_ ) );
BUF_X1 \myifu/_1978_ ( .A(\araddr_IFU [10] ), .Z(\myifu/_0042_ ) );
BUF_X1 \myifu/_1979_ ( .A(\pc_jump [11] ), .Z(\myifu/_0866_ ) );
BUF_X1 \myifu/_1980_ ( .A(\araddr_IFU [11] ), .Z(\myifu/_0043_ ) );
BUF_X1 \myifu/_1981_ ( .A(\pc_jump [12] ), .Z(\myifu/_0867_ ) );
BUF_X1 \myifu/_1982_ ( .A(\araddr_IFU [12] ), .Z(\myifu/_0044_ ) );
BUF_X1 \myifu/_1983_ ( .A(\pc_jump [13] ), .Z(\myifu/_0868_ ) );
BUF_X1 \myifu/_1984_ ( .A(\araddr_IFU [13] ), .Z(\myifu/_0045_ ) );
BUF_X1 \myifu/_1985_ ( .A(\pc_jump [14] ), .Z(\myifu/_0869_ ) );
BUF_X1 \myifu/_1986_ ( .A(\araddr_IFU [14] ), .Z(\myifu/_0046_ ) );
BUF_X1 \myifu/_1987_ ( .A(\pc_jump [15] ), .Z(\myifu/_0870_ ) );
BUF_X1 \myifu/_1988_ ( .A(\araddr_IFU [15] ), .Z(\myifu/_0047_ ) );
BUF_X1 \myifu/_1989_ ( .A(\pc_jump [16] ), .Z(\myifu/_0871_ ) );
BUF_X1 \myifu/_1990_ ( .A(\araddr_IFU [16] ), .Z(\myifu/_0048_ ) );
BUF_X1 \myifu/_1991_ ( .A(\pc_jump [17] ), .Z(\myifu/_0872_ ) );
BUF_X1 \myifu/_1992_ ( .A(\araddr_IFU [17] ), .Z(\myifu/_0049_ ) );
BUF_X1 \myifu/_1993_ ( .A(\pc_jump [18] ), .Z(\myifu/_0873_ ) );
BUF_X1 \myifu/_1994_ ( .A(\araddr_IFU [18] ), .Z(\myifu/_0050_ ) );
BUF_X1 \myifu/_1995_ ( .A(\pc_jump [19] ), .Z(\myifu/_0874_ ) );
BUF_X1 \myifu/_1996_ ( .A(\araddr_IFU [19] ), .Z(\myifu/_0051_ ) );
BUF_X1 \myifu/_1997_ ( .A(\pc_jump [20] ), .Z(\myifu/_0876_ ) );
BUF_X1 \myifu/_1998_ ( .A(\araddr_IFU [20] ), .Z(\myifu/_0052_ ) );
BUF_X1 \myifu/_1999_ ( .A(\pc_jump [21] ), .Z(\myifu/_0877_ ) );
BUF_X1 \myifu/_2000_ ( .A(\araddr_IFU [21] ), .Z(\myifu/_0053_ ) );
BUF_X1 \myifu/_2001_ ( .A(\pc_jump [22] ), .Z(\myifu/_0878_ ) );
BUF_X1 \myifu/_2002_ ( .A(\araddr_IFU [22] ), .Z(\myifu/_0054_ ) );
BUF_X1 \myifu/_2003_ ( .A(\pc_jump [23] ), .Z(\myifu/_0879_ ) );
BUF_X1 \myifu/_2004_ ( .A(\araddr_IFU [23] ), .Z(\myifu/_0055_ ) );
BUF_X1 \myifu/_2005_ ( .A(\pc_jump [24] ), .Z(\myifu/_0880_ ) );
BUF_X1 \myifu/_2006_ ( .A(\araddr_IFU [24] ), .Z(\myifu/_0056_ ) );
BUF_X1 \myifu/_2007_ ( .A(\pc_jump [25] ), .Z(\myifu/_0881_ ) );
BUF_X1 \myifu/_2008_ ( .A(\araddr_IFU [25] ), .Z(\myifu/_0057_ ) );
BUF_X1 \myifu/_2009_ ( .A(\pc_jump [26] ), .Z(\myifu/_0882_ ) );
BUF_X1 \myifu/_2010_ ( .A(\araddr_IFU [26] ), .Z(\myifu/_0058_ ) );
BUF_X1 \myifu/_2011_ ( .A(\pc_jump [27] ), .Z(\myifu/_0883_ ) );
BUF_X1 \myifu/_2012_ ( .A(\araddr_IFU [27] ), .Z(\myifu/_0059_ ) );
BUF_X1 \myifu/_2013_ ( .A(\pc_jump [28] ), .Z(\myifu/_0884_ ) );
BUF_X1 \myifu/_2014_ ( .A(\araddr_IFU [28] ), .Z(\myifu/_0060_ ) );
BUF_X1 \myifu/_2015_ ( .A(\pc_jump [29] ), .Z(\myifu/_0885_ ) );
BUF_X1 \myifu/_2016_ ( .A(\araddr_IFU [29] ), .Z(\myifu/_0061_ ) );
BUF_X1 \myifu/_2017_ ( .A(\pc_jump [30] ), .Z(\myifu/_0887_ ) );
BUF_X1 \myifu/_2018_ ( .A(\araddr_IFU [30] ), .Z(\myifu/_0062_ ) );
BUF_X1 \myifu/_2019_ ( .A(\pc_jump [31] ), .Z(\myifu/_0888_ ) );
BUF_X1 \myifu/_2020_ ( .A(\araddr_IFU [31] ), .Z(\myifu/_0063_ ) );
BUF_X1 \myifu/_2021_ ( .A(check_quest ), .Z(\myifu/_0141_ ) );
BUF_X1 \myifu/_2022_ ( .A(\myifu/state [1] ), .Z(\myifu/_0943_ ) );
BUF_X1 \myifu/_2023_ ( .A(\myifu/_0973_ ), .Z(IFU_valid_IDU ) );
BUF_X1 \myifu/_2024_ ( .A(\myifu/_0025_ ), .Z(\myifu/_0004_ ) );
BUF_X1 \myifu/_2025_ ( .A(\rresp_IFU [1] ), .Z(\myifu/_0939_ ) );
BUF_X1 \myifu/_2026_ ( .A(\rresp_IFU [0] ), .Z(\myifu/_0938_ ) );
BUF_X1 \myifu/_2027_ ( .A(rvalid_IFU ), .Z(\myifu/_0940_ ) );
BUF_X1 \myifu/_2028_ ( .A(rlast_IFU ), .Z(\myifu/_0935_ ) );
BUF_X1 \myifu/_2029_ ( .A(\rid_IFU [1] ), .Z(\myifu/_0932_ ) );
BUF_X1 \myifu/_2030_ ( .A(\rid_IFU [0] ), .Z(\myifu/_0931_ ) );
BUF_X1 \myifu/_2031_ ( .A(\rid_IFU [3] ), .Z(\myifu/_0934_ ) );
BUF_X1 \myifu/_2032_ ( .A(\rid_IFU [2] ), .Z(\myifu/_0933_ ) );
BUF_X1 \myifu/_2033_ ( .A(\myifu/state [2] ), .Z(\myifu/_0944_ ) );
BUF_X1 \myifu/_2034_ ( .A(IDU_ready_IFU ), .Z(\myifu/_0929_ ) );
BUF_X1 \myifu/_2035_ ( .A(\myifu/tag_out [0] ), .Z(\myifu/_0945_ ) );
BUF_X1 \myifu/_2036_ ( .A(\myifu/tag_out [1] ), .Z(\myifu/_0956_ ) );
BUF_X1 \myifu/_2037_ ( .A(\myifu/tag_out [2] ), .Z(\myifu/_0964_ ) );
BUF_X1 \myifu/_2038_ ( .A(\myifu/tag_out [3] ), .Z(\myifu/_0965_ ) );
BUF_X1 \myifu/_2039_ ( .A(\myifu/tag_out [4] ), .Z(\myifu/_0966_ ) );
BUF_X1 \myifu/_2040_ ( .A(\myifu/tag_out [5] ), .Z(\myifu/_0967_ ) );
BUF_X1 \myifu/_2041_ ( .A(\myifu/tag_out [6] ), .Z(\myifu/_0968_ ) );
BUF_X1 \myifu/_2042_ ( .A(\myifu/tag_out [7] ), .Z(\myifu/_0969_ ) );
BUF_X1 \myifu/_2043_ ( .A(\myifu/tag_out [8] ), .Z(\myifu/_0970_ ) );
BUF_X1 \myifu/_2044_ ( .A(\myifu/tag_out [9] ), .Z(\myifu/_0971_ ) );
BUF_X1 \myifu/_2045_ ( .A(\myifu/tag_out [10] ), .Z(\myifu/_0946_ ) );
BUF_X1 \myifu/_2046_ ( .A(\myifu/tag_out [11] ), .Z(\myifu/_0947_ ) );
BUF_X1 \myifu/_2047_ ( .A(\myifu/tag_out [12] ), .Z(\myifu/_0948_ ) );
BUF_X1 \myifu/_2048_ ( .A(\myifu/tag_out [13] ), .Z(\myifu/_0949_ ) );
BUF_X1 \myifu/_2049_ ( .A(\myifu/tag_out [14] ), .Z(\myifu/_0950_ ) );
BUF_X1 \myifu/_2050_ ( .A(\myifu/tag_out [15] ), .Z(\myifu/_0951_ ) );
BUF_X1 \myifu/_2051_ ( .A(\myifu/tag_out [16] ), .Z(\myifu/_0952_ ) );
BUF_X1 \myifu/_2052_ ( .A(\myifu/tag_out [17] ), .Z(\myifu/_0953_ ) );
BUF_X1 \myifu/_2053_ ( .A(\myifu/tag_out [18] ), .Z(\myifu/_0954_ ) );
BUF_X1 \myifu/_2054_ ( .A(\myifu/tag_out [19] ), .Z(\myifu/_0955_ ) );
BUF_X1 \myifu/_2055_ ( .A(\myifu/tag_out [20] ), .Z(\myifu/_0957_ ) );
BUF_X1 \myifu/_2056_ ( .A(\myifu/tag_out [21] ), .Z(\myifu/_0958_ ) );
BUF_X1 \myifu/_2057_ ( .A(\myifu/tag_out [22] ), .Z(\myifu/_0959_ ) );
BUF_X1 \myifu/_2058_ ( .A(\myifu/tag_out [23] ), .Z(\myifu/_0960_ ) );
BUF_X1 \myifu/_2059_ ( .A(\myifu/tag_out [24] ), .Z(\myifu/_0961_ ) );
BUF_X1 \myifu/_2060_ ( .A(\myifu/tag_out [25] ), .Z(\myifu/_0962_ ) );
BUF_X1 \myifu/_2061_ ( .A(\myifu/tag_out [26] ), .Z(\myifu/_0963_ ) );
BUF_X1 \myifu/_2062_ ( .A(\myifu/valid_out ), .Z(\myifu/_0975_ ) );
BUF_X1 \myifu/_2063_ ( .A(\myifu/_0022_ ), .Z(\myifu/_0001_ ) );
BUF_X1 \myifu/_2064_ ( .A(arready_IFU ), .Z(\myifu/_0071_ ) );
BUF_X1 \myifu/_2065_ ( .A(\myifu/_0023_ ), .Z(\myifu/_0002_ ) );
BUF_X1 \myifu/_2066_ ( .A(\myifu/_0021_ ), .Z(\myifu/_0000_ ) );
BUF_X1 \myifu/_2067_ ( .A(\myifu/_0937_ ), .Z(rready_IFU ) );
BUF_X1 \myifu/_2068_ ( .A(\myifu/_0936_ ), .Z(rmem_quest_IFU ) );
BUF_X1 \myifu/_2069_ ( .A(\myifu/valid_in ), .Z(\myifu/_0974_ ) );
BUF_X1 \myifu/_2070_ ( .A(\myifu/_0858_ ), .Z(\myifu/offset [0] ) );
BUF_X1 \myifu/_2071_ ( .A(\myifu/_0859_ ), .Z(\myifu/offset [1] ) );
BUF_X1 \myifu/_2072_ ( .A(\myifu/tmp_offset [2] ), .Z(\myifu/_0972_ ) );
BUF_X1 \myifu/_2073_ ( .A(\myifu/_0860_ ), .Z(\myifu/offset [2] ) );
BUF_X1 \myifu/_2074_ ( .A(\myifu/_0005_ ), .Z(\myifu/_0026_ ) );
BUF_X1 \myifu/_2075_ ( .A(\IF_ID_inst [0] ), .Z(\myifu/_0174_ ) );
BUF_X1 \myifu/_2076_ ( .A(\rdata_IFU [0] ), .Z(\myifu/_0897_ ) );
BUF_X1 \myifu/_2077_ ( .A(\myifu/data_out [0] ), .Z(\myifu/_0142_ ) );
BUF_X1 \myifu/_2078_ ( .A(\IF_ID_inst [1] ), .Z(\myifu/_0185_ ) );
BUF_X1 \myifu/_2079_ ( .A(\rdata_IFU [1] ), .Z(\myifu/_0908_ ) );
BUF_X1 \myifu/_2080_ ( .A(\myifu/data_out [1] ), .Z(\myifu/_0153_ ) );
BUF_X1 \myifu/_2081_ ( .A(\IF_ID_inst [2] ), .Z(\myifu/_0196_ ) );
BUF_X1 \myifu/_2082_ ( .A(\rdata_IFU [2] ), .Z(\myifu/_0919_ ) );
BUF_X1 \myifu/_2083_ ( .A(\myifu/data_out [2] ), .Z(\myifu/_0164_ ) );
BUF_X1 \myifu/_2084_ ( .A(\IF_ID_inst [3] ), .Z(\myifu/_0198_ ) );
BUF_X1 \myifu/_2085_ ( .A(\rdata_IFU [3] ), .Z(\myifu/_0922_ ) );
BUF_X1 \myifu/_2086_ ( .A(\myifu/data_out [3] ), .Z(\myifu/_0167_ ) );
BUF_X1 \myifu/_2087_ ( .A(\IF_ID_inst [4] ), .Z(\myifu/_0199_ ) );
BUF_X1 \myifu/_2088_ ( .A(\rdata_IFU [4] ), .Z(\myifu/_0923_ ) );
BUF_X1 \myifu/_2089_ ( .A(\myifu/data_out [4] ), .Z(\myifu/_0168_ ) );
BUF_X1 \myifu/_2090_ ( .A(\IF_ID_inst [5] ), .Z(\myifu/_0200_ ) );
BUF_X1 \myifu/_2091_ ( .A(\rdata_IFU [5] ), .Z(\myifu/_0924_ ) );
BUF_X1 \myifu/_2092_ ( .A(\myifu/data_out [5] ), .Z(\myifu/_0169_ ) );
BUF_X1 \myifu/_2093_ ( .A(\IF_ID_inst [6] ), .Z(\myifu/_0201_ ) );
BUF_X1 \myifu/_2094_ ( .A(\rdata_IFU [6] ), .Z(\myifu/_0925_ ) );
BUF_X1 \myifu/_2095_ ( .A(\myifu/data_out [6] ), .Z(\myifu/_0170_ ) );
BUF_X1 \myifu/_2096_ ( .A(\IF_ID_inst [7] ), .Z(\myifu/_0202_ ) );
BUF_X1 \myifu/_2097_ ( .A(\rdata_IFU [7] ), .Z(\myifu/_0926_ ) );
BUF_X1 \myifu/_2098_ ( .A(\myifu/data_out [7] ), .Z(\myifu/_0171_ ) );
BUF_X1 \myifu/_2099_ ( .A(\IF_ID_inst [8] ), .Z(\myifu/_0203_ ) );
BUF_X1 \myifu/_2100_ ( .A(\rdata_IFU [8] ), .Z(\myifu/_0927_ ) );
BUF_X1 \myifu/_2101_ ( .A(\myifu/data_out [8] ), .Z(\myifu/_0172_ ) );
BUF_X1 \myifu/_2102_ ( .A(\IF_ID_inst [9] ), .Z(\myifu/_0204_ ) );
BUF_X1 \myifu/_2103_ ( .A(\rdata_IFU [9] ), .Z(\myifu/_0928_ ) );
BUF_X1 \myifu/_2104_ ( .A(\myifu/data_out [9] ), .Z(\myifu/_0173_ ) );
BUF_X1 \myifu/_2105_ ( .A(\IF_ID_inst [10] ), .Z(\myifu/_0175_ ) );
BUF_X1 \myifu/_2106_ ( .A(\rdata_IFU [10] ), .Z(\myifu/_0898_ ) );
BUF_X1 \myifu/_2107_ ( .A(\myifu/data_out [10] ), .Z(\myifu/_0143_ ) );
BUF_X1 \myifu/_2108_ ( .A(\IF_ID_inst [11] ), .Z(\myifu/_0176_ ) );
BUF_X1 \myifu/_2109_ ( .A(\rdata_IFU [11] ), .Z(\myifu/_0899_ ) );
BUF_X1 \myifu/_2110_ ( .A(\myifu/data_out [11] ), .Z(\myifu/_0144_ ) );
BUF_X1 \myifu/_2111_ ( .A(\IF_ID_inst [12] ), .Z(\myifu/_0177_ ) );
BUF_X1 \myifu/_2112_ ( .A(\rdata_IFU [12] ), .Z(\myifu/_0900_ ) );
BUF_X1 \myifu/_2113_ ( .A(\myifu/data_out [12] ), .Z(\myifu/_0145_ ) );
BUF_X1 \myifu/_2114_ ( .A(\IF_ID_inst [13] ), .Z(\myifu/_0178_ ) );
BUF_X1 \myifu/_2115_ ( .A(\rdata_IFU [13] ), .Z(\myifu/_0901_ ) );
BUF_X1 \myifu/_2116_ ( .A(\myifu/data_out [13] ), .Z(\myifu/_0146_ ) );
BUF_X1 \myifu/_2117_ ( .A(\IF_ID_inst [14] ), .Z(\myifu/_0179_ ) );
BUF_X1 \myifu/_2118_ ( .A(\rdata_IFU [14] ), .Z(\myifu/_0902_ ) );
BUF_X1 \myifu/_2119_ ( .A(\myifu/data_out [14] ), .Z(\myifu/_0147_ ) );
BUF_X1 \myifu/_2120_ ( .A(\IF_ID_inst [15] ), .Z(\myifu/_0180_ ) );
BUF_X1 \myifu/_2121_ ( .A(\rdata_IFU [15] ), .Z(\myifu/_0903_ ) );
BUF_X1 \myifu/_2122_ ( .A(\myifu/data_out [15] ), .Z(\myifu/_0148_ ) );
BUF_X1 \myifu/_2123_ ( .A(\IF_ID_inst [16] ), .Z(\myifu/_0181_ ) );
BUF_X1 \myifu/_2124_ ( .A(\rdata_IFU [16] ), .Z(\myifu/_0904_ ) );
BUF_X1 \myifu/_2125_ ( .A(\myifu/data_out [16] ), .Z(\myifu/_0149_ ) );
BUF_X1 \myifu/_2126_ ( .A(\IF_ID_inst [17] ), .Z(\myifu/_0182_ ) );
BUF_X1 \myifu/_2127_ ( .A(\rdata_IFU [17] ), .Z(\myifu/_0905_ ) );
BUF_X1 \myifu/_2128_ ( .A(\myifu/data_out [17] ), .Z(\myifu/_0150_ ) );
BUF_X1 \myifu/_2129_ ( .A(\IF_ID_inst [18] ), .Z(\myifu/_0183_ ) );
BUF_X1 \myifu/_2130_ ( .A(\rdata_IFU [18] ), .Z(\myifu/_0906_ ) );
BUF_X1 \myifu/_2131_ ( .A(\myifu/data_out [18] ), .Z(\myifu/_0151_ ) );
BUF_X1 \myifu/_2132_ ( .A(\IF_ID_inst [19] ), .Z(\myifu/_0184_ ) );
BUF_X1 \myifu/_2133_ ( .A(\rdata_IFU [19] ), .Z(\myifu/_0907_ ) );
BUF_X1 \myifu/_2134_ ( .A(\myifu/data_out [19] ), .Z(\myifu/_0152_ ) );
BUF_X1 \myifu/_2135_ ( .A(\IF_ID_inst [20] ), .Z(\myifu/_0186_ ) );
BUF_X1 \myifu/_2136_ ( .A(\rdata_IFU [20] ), .Z(\myifu/_0909_ ) );
BUF_X1 \myifu/_2137_ ( .A(\myifu/data_out [20] ), .Z(\myifu/_0154_ ) );
BUF_X1 \myifu/_2138_ ( .A(\IF_ID_inst [21] ), .Z(\myifu/_0187_ ) );
BUF_X1 \myifu/_2139_ ( .A(\rdata_IFU [21] ), .Z(\myifu/_0910_ ) );
BUF_X1 \myifu/_2140_ ( .A(\myifu/data_out [21] ), .Z(\myifu/_0155_ ) );
BUF_X1 \myifu/_2141_ ( .A(\IF_ID_inst [22] ), .Z(\myifu/_0188_ ) );
BUF_X1 \myifu/_2142_ ( .A(\rdata_IFU [22] ), .Z(\myifu/_0911_ ) );
BUF_X1 \myifu/_2143_ ( .A(\myifu/data_out [22] ), .Z(\myifu/_0156_ ) );
BUF_X1 \myifu/_2144_ ( .A(\IF_ID_inst [23] ), .Z(\myifu/_0189_ ) );
BUF_X1 \myifu/_2145_ ( .A(\rdata_IFU [23] ), .Z(\myifu/_0912_ ) );
BUF_X1 \myifu/_2146_ ( .A(\myifu/data_out [23] ), .Z(\myifu/_0157_ ) );
BUF_X1 \myifu/_2147_ ( .A(\IF_ID_inst [24] ), .Z(\myifu/_0190_ ) );
BUF_X1 \myifu/_2148_ ( .A(\rdata_IFU [24] ), .Z(\myifu/_0913_ ) );
BUF_X1 \myifu/_2149_ ( .A(\myifu/data_out [24] ), .Z(\myifu/_0158_ ) );
BUF_X1 \myifu/_2150_ ( .A(\IF_ID_inst [25] ), .Z(\myifu/_0191_ ) );
BUF_X1 \myifu/_2151_ ( .A(\rdata_IFU [25] ), .Z(\myifu/_0914_ ) );
BUF_X1 \myifu/_2152_ ( .A(\myifu/data_out [25] ), .Z(\myifu/_0159_ ) );
BUF_X1 \myifu/_2153_ ( .A(\IF_ID_inst [26] ), .Z(\myifu/_0192_ ) );
BUF_X1 \myifu/_2154_ ( .A(\rdata_IFU [26] ), .Z(\myifu/_0915_ ) );
BUF_X1 \myifu/_2155_ ( .A(\myifu/data_out [26] ), .Z(\myifu/_0160_ ) );
BUF_X1 \myifu/_2156_ ( .A(\IF_ID_inst [27] ), .Z(\myifu/_0193_ ) );
BUF_X1 \myifu/_2157_ ( .A(\rdata_IFU [27] ), .Z(\myifu/_0916_ ) );
BUF_X1 \myifu/_2158_ ( .A(\myifu/data_out [27] ), .Z(\myifu/_0161_ ) );
BUF_X1 \myifu/_2159_ ( .A(\IF_ID_inst [28] ), .Z(\myifu/_0194_ ) );
BUF_X1 \myifu/_2160_ ( .A(\rdata_IFU [28] ), .Z(\myifu/_0917_ ) );
BUF_X1 \myifu/_2161_ ( .A(\myifu/data_out [28] ), .Z(\myifu/_0162_ ) );
BUF_X1 \myifu/_2162_ ( .A(\IF_ID_inst [29] ), .Z(\myifu/_0195_ ) );
BUF_X1 \myifu/_2163_ ( .A(\rdata_IFU [29] ), .Z(\myifu/_0918_ ) );
BUF_X1 \myifu/_2164_ ( .A(\myifu/data_out [29] ), .Z(\myifu/_0163_ ) );
BUF_X1 \myifu/_2165_ ( .A(\IF_ID_inst [30] ), .Z(\myifu/_0197_ ) );
BUF_X1 \myifu/_2166_ ( .A(\rdata_IFU [30] ), .Z(\myifu/_0920_ ) );
BUF_X1 \myifu/_2167_ ( .A(\myifu/data_out [30] ), .Z(\myifu/_0165_ ) );
BUF_X1 \myifu/_2168_ ( .A(\myifu/pred_jump ), .Z(\myifu/_0896_ ) );
BUF_X1 \myifu/_2169_ ( .A(\rdata_IFU [31] ), .Z(\myifu/_0921_ ) );
BUF_X1 \myifu/_2170_ ( .A(\myifu/data_out [31] ), .Z(\myifu/_0166_ ) );
BUF_X1 \myifu/_2171_ ( .A(\myifu/_0007_ ), .Z(\myifu/_0028_ ) );
BUF_X1 \myifu/_2172_ ( .A(\myifu/_0006_ ), .Z(\myifu/_0027_ ) );
BUF_X1 \myifu/_2173_ ( .A(\myifu/_0008_ ), .Z(\myifu/_0029_ ) );
BUF_X1 \myifu/_2174_ ( .A(\myifu/_0009_ ), .Z(\myifu/_0030_ ) );
BUF_X1 \myifu/_2175_ ( .A(\myifu/_0010_ ), .Z(\myifu/_0031_ ) );
BUF_X1 \myifu/_2176_ ( .A(\myifu/_0011_ ), .Z(\myifu/_0032_ ) );
BUF_X1 \myifu/_2177_ ( .A(\myifu/_0012_ ), .Z(\myifu/_0033_ ) );
BUF_X1 \myifu/_2178_ ( .A(\myifu/_0013_ ), .Z(\myifu/_0034_ ) );
BUF_X1 \myifu/_2179_ ( .A(\myifu/_0014_ ), .Z(\myifu/_0035_ ) );
BUF_X1 \myifu/_2180_ ( .A(\myifu/_0015_ ), .Z(\myifu/_0036_ ) );
BUF_X1 \myifu/_2181_ ( .A(\myifu/_0016_ ), .Z(\myifu/_0037_ ) );
BUF_X1 \myifu/_2182_ ( .A(\myifu/_0017_ ), .Z(\myifu/_0038_ ) );
BUF_X1 \myifu/_2183_ ( .A(\myifu/_0018_ ), .Z(\myifu/_0039_ ) );
BUF_X1 \myifu/_2184_ ( .A(\myifu/_0019_ ), .Z(\myifu/_0040_ ) );
BUF_X1 \myifu/_2185_ ( .A(\myifu/_0020_ ), .Z(\myifu/_0041_ ) );
BUF_X1 \myifu/_2186_ ( .A(\myifu/_0106_ ), .Z(\myifu/_1064_ ) );
BUF_X1 \myifu/_2187_ ( .A(\myifu/_0107_ ), .Z(\myifu/_1065_ ) );
BUF_X1 \myifu/_2188_ ( .A(\myifu/_0108_ ), .Z(\myifu/_1066_ ) );
BUF_X1 \myifu/_2189_ ( .A(\myifu/_0109_ ), .Z(\myifu/_1067_ ) );
BUF_X1 \myifu/_2190_ ( .A(\myifu/_0110_ ), .Z(\myifu/_1068_ ) );
BUF_X1 \myifu/_2191_ ( .A(\myifu/_0111_ ), .Z(\myifu/_1069_ ) );
BUF_X1 \myifu/_2192_ ( .A(\myifu/_0112_ ), .Z(\myifu/_1070_ ) );
BUF_X1 \myifu/_2193_ ( .A(\myifu/_0113_ ), .Z(\myifu/_1071_ ) );
BUF_X1 \myifu/_2194_ ( .A(\myifu/_0114_ ), .Z(\myifu/_1072_ ) );
BUF_X1 \myifu/_2195_ ( .A(\myifu/_0115_ ), .Z(\myifu/_1073_ ) );
BUF_X1 \myifu/_2196_ ( .A(\myifu/_0116_ ), .Z(\myifu/_1074_ ) );
BUF_X1 \myifu/_2197_ ( .A(\myifu/_0117_ ), .Z(\myifu/_1075_ ) );
BUF_X1 \myifu/_2198_ ( .A(\myifu/_0118_ ), .Z(\myifu/_1076_ ) );
BUF_X1 \myifu/_2199_ ( .A(\myifu/_0119_ ), .Z(\myifu/_1077_ ) );
BUF_X1 \myifu/_2200_ ( .A(\myifu/_0120_ ), .Z(\myifu/_1078_ ) );
BUF_X1 \myifu/_2201_ ( .A(\myifu/_0121_ ), .Z(\myifu/_1079_ ) );
BUF_X1 \myifu/_2202_ ( .A(\myifu/_0122_ ), .Z(\myifu/_1080_ ) );
BUF_X1 \myifu/_2203_ ( .A(\myifu/_0123_ ), .Z(\myifu/_1081_ ) );
BUF_X1 \myifu/_2204_ ( .A(\myifu/_0124_ ), .Z(\myifu/_1082_ ) );
BUF_X1 \myifu/_2205_ ( .A(\myifu/_0125_ ), .Z(\myifu/_1083_ ) );
BUF_X1 \myifu/_2206_ ( .A(\myifu/_0126_ ), .Z(\myifu/_1084_ ) );
BUF_X1 \myifu/_2207_ ( .A(\myifu/_0127_ ), .Z(\myifu/_1085_ ) );
BUF_X1 \myifu/_2208_ ( .A(\myifu/_0128_ ), .Z(\myifu/_1086_ ) );
BUF_X1 \myifu/_2209_ ( .A(\myifu/_0129_ ), .Z(\myifu/_1087_ ) );
BUF_X1 \myifu/_2210_ ( .A(\myifu/_0130_ ), .Z(\myifu/_1088_ ) );
BUF_X1 \myifu/_2211_ ( .A(\myifu/_0131_ ), .Z(\myifu/_1089_ ) );
BUF_X1 \myifu/_2212_ ( .A(\myifu/_0132_ ), .Z(\myifu/_1090_ ) );
BUF_X1 \myifu/_2213_ ( .A(\myifu/_0133_ ), .Z(\myifu/_1091_ ) );
BUF_X1 \myifu/_2214_ ( .A(\myifu/_0134_ ), .Z(\myifu/_1092_ ) );
BUF_X1 \myifu/_2215_ ( .A(\myifu/_0135_ ), .Z(\myifu/_1093_ ) );
BUF_X1 \myifu/_2216_ ( .A(\myifu/_0136_ ), .Z(\myifu/_1094_ ) );
BUF_X1 \myifu/_2217_ ( .A(\myifu/_0137_ ), .Z(\myifu/_1095_ ) );
BUF_X1 \myifu/_2218_ ( .A(\myifu/_0003_ ), .Z(\myifu/_0024_ ) );
BUF_X1 \myifu/_2219_ ( .A(check_assert ), .Z(\myifu/_0140_ ) );
BUF_X1 \myifu/_2220_ ( .A(\myifu/_0139_ ), .Z(\myifu/_1097_ ) );
BUF_X1 \myifu/_2221_ ( .A(\myifu/_0073_ ), .Z(\myifu/_1031_ ) );
BUF_X1 \myifu/_2222_ ( .A(\myifu/_0074_ ), .Z(\myifu/_1032_ ) );
BUF_X1 \myifu/_2223_ ( .A(\myifu/_0075_ ), .Z(\myifu/_1033_ ) );
BUF_X1 \myifu/_2224_ ( .A(\myifu/_0076_ ), .Z(\myifu/_1034_ ) );
BUF_X1 \myifu/_2225_ ( .A(\myifu/_0077_ ), .Z(\myifu/_1035_ ) );
BUF_X1 \myifu/_2226_ ( .A(\myifu/_0078_ ), .Z(\myifu/_1036_ ) );
BUF_X1 \myifu/_2227_ ( .A(\myifu/_0079_ ), .Z(\myifu/_1037_ ) );
BUF_X1 \myifu/_2228_ ( .A(\myifu/_0080_ ), .Z(\myifu/_1038_ ) );
BUF_X1 \myifu/_2229_ ( .A(\myifu/_0081_ ), .Z(\myifu/_1039_ ) );
BUF_X1 \myifu/_2230_ ( .A(\myifu/_0082_ ), .Z(\myifu/_1040_ ) );
BUF_X1 \myifu/_2231_ ( .A(\myifu/_0083_ ), .Z(\myifu/_1041_ ) );
BUF_X1 \myifu/_2232_ ( .A(\myifu/_0084_ ), .Z(\myifu/_1042_ ) );
BUF_X1 \myifu/_2233_ ( .A(\myifu/_0085_ ), .Z(\myifu/_1043_ ) );
BUF_X1 \myifu/_2234_ ( .A(\myifu/_0086_ ), .Z(\myifu/_1044_ ) );
BUF_X1 \myifu/_2235_ ( .A(\myifu/_0087_ ), .Z(\myifu/_1045_ ) );
BUF_X1 \myifu/_2236_ ( .A(\myifu/_0088_ ), .Z(\myifu/_1046_ ) );
BUF_X1 \myifu/_2237_ ( .A(\myifu/_0089_ ), .Z(\myifu/_1047_ ) );
BUF_X1 \myifu/_2238_ ( .A(\myifu/_0090_ ), .Z(\myifu/_1048_ ) );
BUF_X1 \myifu/_2239_ ( .A(\myifu/_0091_ ), .Z(\myifu/_1049_ ) );
BUF_X1 \myifu/_2240_ ( .A(\myifu/_0092_ ), .Z(\myifu/_1050_ ) );
BUF_X1 \myifu/_2241_ ( .A(\myifu/_0093_ ), .Z(\myifu/_1051_ ) );
BUF_X1 \myifu/_2242_ ( .A(\myifu/_0094_ ), .Z(\myifu/_1052_ ) );
BUF_X1 \myifu/_2243_ ( .A(\myifu/_0095_ ), .Z(\myifu/_1053_ ) );
BUF_X1 \myifu/_2244_ ( .A(\myifu/_0096_ ), .Z(\myifu/_1054_ ) );
BUF_X1 \myifu/_2245_ ( .A(\myifu/_0097_ ), .Z(\myifu/_1055_ ) );
BUF_X1 \myifu/_2246_ ( .A(\myifu/_0098_ ), .Z(\myifu/_1056_ ) );
BUF_X1 \myifu/_2247_ ( .A(\myifu/_0099_ ), .Z(\myifu/_1057_ ) );
BUF_X1 \myifu/_2248_ ( .A(\myifu/_0100_ ), .Z(\myifu/_1058_ ) );
BUF_X1 \myifu/_2249_ ( .A(\myifu/_0101_ ), .Z(\myifu/_1059_ ) );
BUF_X1 \myifu/_2250_ ( .A(\myifu/_0102_ ), .Z(\myifu/_1060_ ) );
BUF_X1 \myifu/_2251_ ( .A(\myifu/_0103_ ), .Z(\myifu/_1061_ ) );
BUF_X1 \myifu/_2252_ ( .A(\myifu/_0104_ ), .Z(\myifu/_1062_ ) );
BUF_X1 \myifu/_2253_ ( .A(\myifu/_0105_ ), .Z(\myifu/_1063_ ) );
BUF_X1 \myifu/_2254_ ( .A(\myifu/_0138_ ), .Z(\myifu/_1096_ ) );
INV_X32 \myifu/myicache/_1970_ ( .A(\myifu/myicache/_0689_ ), .ZN(\myifu/myicache/_0956_ ) );
AND2_X4 \myifu/myicache/_1971_ ( .A1(\myifu/myicache/_0956_ ), .A2(fanout_net_20 ), .ZN(\myifu/myicache/_0957_ ) );
BUF_X4 \myifu/myicache/_1972_ ( .A(\myifu/myicache/_0957_ ), .Z(\myifu/myicache/_0958_ ) );
BUF_X4 \myifu/myicache/_1973_ ( .A(\myifu/myicache/_0958_ ), .Z(\myifu/myicache/_0959_ ) );
NOR2_X4 \myifu/myicache/_1974_ ( .A1(\myifu/myicache/_0956_ ), .A2(fanout_net_20 ), .ZN(\myifu/myicache/_0960_ ) );
BUF_X4 \myifu/myicache/_1975_ ( .A(\myifu/myicache/_0960_ ), .Z(\myifu/myicache/_0961_ ) );
AOI22_X1 \myifu/myicache/_1976_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1092_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1119_ ), .ZN(\myifu/myicache/_0962_ ) );
NOR2_X4 \myifu/myicache/_1977_ ( .A1(fanout_net_20 ), .A2(\myifu/myicache/_0689_ ), .ZN(\myifu/myicache/_0963_ ) );
BUF_X4 \myifu/myicache/_1978_ ( .A(\myifu/myicache/_0963_ ), .Z(\myifu/myicache/_0964_ ) );
NAND2_X1 \myifu/myicache/_1979_ ( .A1(\myifu/myicache/_0964_ ), .A2(\myifu/myicache/_1065_ ), .ZN(\myifu/myicache/_0965_ ) );
NAND3_X1 \myifu/myicache/_1980_ ( .A1(fanout_net_20 ), .A2(\myifu/myicache/_0689_ ), .A3(\myifu/myicache/_1146_ ), .ZN(\myifu/myicache/_0966_ ) );
NAND3_X1 \myifu/myicache/_1981_ ( .A1(\myifu/myicache/_0962_ ), .A2(\myifu/myicache/_0965_ ), .A3(\myifu/myicache/_0966_ ), .ZN(\myifu/myicache/_1200_ ) );
BUF_X4 \myifu/myicache/_1982_ ( .A(\myifu/myicache/_0958_ ), .Z(\myifu/myicache/_0967_ ) );
BUF_X4 \myifu/myicache/_1983_ ( .A(\myifu/myicache/_0960_ ), .Z(\myifu/myicache/_0968_ ) );
AOI22_X1 \myifu/myicache/_1984_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1103_ ), .B1(\myifu/myicache/_0968_ ), .B2(\myifu/myicache/_1130_ ), .ZN(\myifu/myicache/_0969_ ) );
AND2_X4 \myifu/myicache/_1985_ ( .A1(fanout_net_20 ), .A2(\myifu/myicache/_0689_ ), .ZN(\myifu/myicache/_0970_ ) );
BUF_X8 \myifu/myicache/_1986_ ( .A(\myifu/myicache/_0970_ ), .Z(\myifu/myicache/_0971_ ) );
BUF_X4 \myifu/myicache/_1987_ ( .A(\myifu/myicache/_0971_ ), .Z(\myifu/myicache/_0972_ ) );
AOI22_X1 \myifu/myicache/_1988_ ( .A1(\myifu/myicache/_1157_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1076_ ), .ZN(\myifu/myicache/_0973_ ) );
NAND2_X1 \myifu/myicache/_1989_ ( .A1(\myifu/myicache/_0969_ ), .A2(\myifu/myicache/_0973_ ), .ZN(\myifu/myicache/_1211_ ) );
BUF_X4 \myifu/myicache/_1990_ ( .A(\myifu/myicache/_0971_ ), .Z(\myifu/myicache/_0974_ ) );
AOI22_X1 \myifu/myicache/_1991_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1111_ ), .B1(\myifu/myicache/_1165_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_0975_ ) );
AOI22_X1 \myifu/myicache/_1992_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1138_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1084_ ), .ZN(\myifu/myicache/_0976_ ) );
NAND2_X1 \myifu/myicache/_1993_ ( .A1(\myifu/myicache/_0975_ ), .A2(\myifu/myicache/_0976_ ), .ZN(\myifu/myicache/_1219_ ) );
AOI22_X1 \myifu/myicache/_1994_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1112_ ), .B1(\myifu/myicache/_1166_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_0977_ ) );
AOI22_X1 \myifu/myicache/_1995_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1139_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1085_ ), .ZN(\myifu/myicache/_0978_ ) );
NAND2_X1 \myifu/myicache/_1996_ ( .A1(\myifu/myicache/_0977_ ), .A2(\myifu/myicache/_0978_ ), .ZN(\myifu/myicache/_1220_ ) );
AOI22_X1 \myifu/myicache/_1997_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1113_ ), .B1(\myifu/myicache/_0968_ ), .B2(\myifu/myicache/_1140_ ), .ZN(\myifu/myicache/_0979_ ) );
AOI22_X1 \myifu/myicache/_1998_ ( .A1(\myifu/myicache/_1167_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1086_ ), .ZN(\myifu/myicache/_0980_ ) );
NAND2_X1 \myifu/myicache/_1999_ ( .A1(\myifu/myicache/_0979_ ), .A2(\myifu/myicache/_0980_ ), .ZN(\myifu/myicache/_1221_ ) );
BUF_X4 \myifu/myicache/_2000_ ( .A(\myifu/myicache/_0960_ ), .Z(\myifu/myicache/_0981_ ) );
AOI22_X1 \myifu/myicache/_2001_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1114_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1141_ ), .ZN(\myifu/myicache/_0982_ ) );
AOI22_X1 \myifu/myicache/_2002_ ( .A1(\myifu/myicache/_1168_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1087_ ), .ZN(\myifu/myicache/_0983_ ) );
NAND2_X1 \myifu/myicache/_2003_ ( .A1(\myifu/myicache/_0982_ ), .A2(\myifu/myicache/_0983_ ), .ZN(\myifu/myicache/_1222_ ) );
AOI22_X1 \myifu/myicache/_2004_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1115_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1142_ ), .ZN(\myifu/myicache/_0984_ ) );
AOI22_X1 \myifu/myicache/_2005_ ( .A1(\myifu/myicache/_1169_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1088_ ), .ZN(\myifu/myicache/_0985_ ) );
NAND2_X1 \myifu/myicache/_2006_ ( .A1(\myifu/myicache/_0984_ ), .A2(\myifu/myicache/_0985_ ), .ZN(\myifu/myicache/_1223_ ) );
AOI22_X1 \myifu/myicache/_2007_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1116_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1143_ ), .ZN(\myifu/myicache/_0986_ ) );
AOI22_X1 \myifu/myicache/_2008_ ( .A1(\myifu/myicache/_1170_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1089_ ), .ZN(\myifu/myicache/_0987_ ) );
NAND2_X1 \myifu/myicache/_2009_ ( .A1(\myifu/myicache/_0986_ ), .A2(\myifu/myicache/_0987_ ), .ZN(\myifu/myicache/_1224_ ) );
AOI22_X1 \myifu/myicache/_2010_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1117_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1144_ ), .ZN(\myifu/myicache/_0988_ ) );
AOI22_X1 \myifu/myicache/_2011_ ( .A1(\myifu/myicache/_1171_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1090_ ), .ZN(\myifu/myicache/_0989_ ) );
NAND2_X1 \myifu/myicache/_2012_ ( .A1(\myifu/myicache/_0988_ ), .A2(\myifu/myicache/_0989_ ), .ZN(\myifu/myicache/_1225_ ) );
AOI22_X1 \myifu/myicache/_2013_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1118_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1145_ ), .ZN(\myifu/myicache/_0990_ ) );
AOI22_X1 \myifu/myicache/_2014_ ( .A1(\myifu/myicache/_1172_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0964_ ), .B2(\myifu/myicache/_1091_ ), .ZN(\myifu/myicache/_0991_ ) );
NAND2_X1 \myifu/myicache/_2015_ ( .A1(\myifu/myicache/_0990_ ), .A2(\myifu/myicache/_0991_ ), .ZN(\myifu/myicache/_1226_ ) );
AOI22_X1 \myifu/myicache/_2016_ ( .A1(\myifu/myicache/_0967_ ), .A2(\myifu/myicache/_1093_ ), .B1(\myifu/myicache/_1147_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_0992_ ) );
BUF_X4 \myifu/myicache/_2017_ ( .A(\myifu/myicache/_0963_ ), .Z(\myifu/myicache/_0993_ ) );
AOI22_X1 \myifu/myicache/_2018_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1120_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1066_ ), .ZN(\myifu/myicache/_0994_ ) );
NAND2_X1 \myifu/myicache/_2019_ ( .A1(\myifu/myicache/_0992_ ), .A2(\myifu/myicache/_0994_ ), .ZN(\myifu/myicache/_1201_ ) );
BUF_X4 \myifu/myicache/_2020_ ( .A(\myifu/myicache/_0958_ ), .Z(\myifu/myicache/_0995_ ) );
AOI22_X1 \myifu/myicache/_2021_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1094_ ), .B1(\myifu/myicache/_1148_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_0996_ ) );
AOI22_X1 \myifu/myicache/_2022_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1121_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1067_ ), .ZN(\myifu/myicache/_0997_ ) );
NAND2_X1 \myifu/myicache/_2023_ ( .A1(\myifu/myicache/_0996_ ), .A2(\myifu/myicache/_0997_ ), .ZN(\myifu/myicache/_1202_ ) );
AOI22_X1 \myifu/myicache/_2024_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1095_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1122_ ), .ZN(\myifu/myicache/_0998_ ) );
AOI22_X1 \myifu/myicache/_2025_ ( .A1(\myifu/myicache/_1149_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1068_ ), .ZN(\myifu/myicache/_0999_ ) );
NAND2_X1 \myifu/myicache/_2026_ ( .A1(\myifu/myicache/_0998_ ), .A2(\myifu/myicache/_0999_ ), .ZN(\myifu/myicache/_1203_ ) );
AOI22_X1 \myifu/myicache/_2027_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1096_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1123_ ), .ZN(\myifu/myicache/_1000_ ) );
AOI22_X1 \myifu/myicache/_2028_ ( .A1(\myifu/myicache/_1150_ ), .A2(\myifu/myicache/_0972_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1069_ ), .ZN(\myifu/myicache/_1001_ ) );
NAND2_X1 \myifu/myicache/_2029_ ( .A1(\myifu/myicache/_1000_ ), .A2(\myifu/myicache/_1001_ ), .ZN(\myifu/myicache/_1204_ ) );
AOI22_X1 \myifu/myicache/_2030_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1097_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1124_ ), .ZN(\myifu/myicache/_1002_ ) );
BUF_X4 \myifu/myicache/_2031_ ( .A(\myifu/myicache/_0971_ ), .Z(\myifu/myicache/_1003_ ) );
AOI22_X1 \myifu/myicache/_2032_ ( .A1(\myifu/myicache/_1151_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1070_ ), .ZN(\myifu/myicache/_1004_ ) );
NAND2_X1 \myifu/myicache/_2033_ ( .A1(\myifu/myicache/_1002_ ), .A2(\myifu/myicache/_1004_ ), .ZN(\myifu/myicache/_1205_ ) );
AOI22_X1 \myifu/myicache/_2034_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1098_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1125_ ), .ZN(\myifu/myicache/_1005_ ) );
AOI22_X1 \myifu/myicache/_2035_ ( .A1(\myifu/myicache/_1152_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1071_ ), .ZN(\myifu/myicache/_1006_ ) );
NAND2_X1 \myifu/myicache/_2036_ ( .A1(\myifu/myicache/_1005_ ), .A2(\myifu/myicache/_1006_ ), .ZN(\myifu/myicache/_1206_ ) );
AOI22_X1 \myifu/myicache/_2037_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1099_ ), .B1(\myifu/myicache/_0981_ ), .B2(\myifu/myicache/_1126_ ), .ZN(\myifu/myicache/_1007_ ) );
AOI22_X1 \myifu/myicache/_2038_ ( .A1(\myifu/myicache/_1153_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1072_ ), .ZN(\myifu/myicache/_1008_ ) );
NAND2_X1 \myifu/myicache/_2039_ ( .A1(\myifu/myicache/_1007_ ), .A2(\myifu/myicache/_1008_ ), .ZN(\myifu/myicache/_1207_ ) );
AOI22_X1 \myifu/myicache/_2040_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1100_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1127_ ), .ZN(\myifu/myicache/_1009_ ) );
AOI22_X1 \myifu/myicache/_2041_ ( .A1(\myifu/myicache/_1154_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1073_ ), .ZN(\myifu/myicache/_1010_ ) );
NAND2_X1 \myifu/myicache/_2042_ ( .A1(\myifu/myicache/_1009_ ), .A2(\myifu/myicache/_1010_ ), .ZN(\myifu/myicache/_1208_ ) );
AOI22_X1 \myifu/myicache/_2043_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1101_ ), .B1(\myifu/myicache/_1155_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_1011_ ) );
AOI22_X1 \myifu/myicache/_2044_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1128_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1074_ ), .ZN(\myifu/myicache/_1012_ ) );
NAND2_X1 \myifu/myicache/_2045_ ( .A1(\myifu/myicache/_1011_ ), .A2(\myifu/myicache/_1012_ ), .ZN(\myifu/myicache/_1209_ ) );
AOI22_X1 \myifu/myicache/_2046_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1102_ ), .B1(\myifu/myicache/_1156_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_1013_ ) );
AOI22_X1 \myifu/myicache/_2047_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1129_ ), .B1(\myifu/myicache/_0993_ ), .B2(\myifu/myicache/_1075_ ), .ZN(\myifu/myicache/_1014_ ) );
NAND2_X1 \myifu/myicache/_2048_ ( .A1(\myifu/myicache/_1013_ ), .A2(\myifu/myicache/_1014_ ), .ZN(\myifu/myicache/_1210_ ) );
AOI22_X1 \myifu/myicache/_2049_ ( .A1(\myifu/myicache/_0995_ ), .A2(\myifu/myicache/_1104_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1131_ ), .ZN(\myifu/myicache/_1015_ ) );
BUF_X4 \myifu/myicache/_2050_ ( .A(\myifu/myicache/_0963_ ), .Z(\myifu/myicache/_1016_ ) );
AOI22_X1 \myifu/myicache/_2051_ ( .A1(\myifu/myicache/_1158_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1077_ ), .ZN(\myifu/myicache/_1017_ ) );
NAND2_X1 \myifu/myicache/_2052_ ( .A1(\myifu/myicache/_1015_ ), .A2(\myifu/myicache/_1017_ ), .ZN(\myifu/myicache/_1212_ ) );
AOI22_X1 \myifu/myicache/_2053_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1105_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1132_ ), .ZN(\myifu/myicache/_1018_ ) );
AOI22_X1 \myifu/myicache/_2054_ ( .A1(\myifu/myicache/_1159_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1078_ ), .ZN(\myifu/myicache/_1019_ ) );
NAND2_X1 \myifu/myicache/_2055_ ( .A1(\myifu/myicache/_1018_ ), .A2(\myifu/myicache/_1019_ ), .ZN(\myifu/myicache/_1213_ ) );
AOI22_X1 \myifu/myicache/_2056_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1106_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1133_ ), .ZN(\myifu/myicache/_1020_ ) );
AOI22_X1 \myifu/myicache/_2057_ ( .A1(\myifu/myicache/_1160_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1079_ ), .ZN(\myifu/myicache/_1021_ ) );
NAND2_X1 \myifu/myicache/_2058_ ( .A1(\myifu/myicache/_1020_ ), .A2(\myifu/myicache/_1021_ ), .ZN(\myifu/myicache/_1214_ ) );
AOI22_X1 \myifu/myicache/_2059_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1107_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1134_ ), .ZN(\myifu/myicache/_1022_ ) );
AOI22_X1 \myifu/myicache/_2060_ ( .A1(\myifu/myicache/_1161_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1080_ ), .ZN(\myifu/myicache/_1023_ ) );
NAND2_X1 \myifu/myicache/_2061_ ( .A1(\myifu/myicache/_1022_ ), .A2(\myifu/myicache/_1023_ ), .ZN(\myifu/myicache/_1215_ ) );
AOI22_X1 \myifu/myicache/_2062_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1108_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1135_ ), .ZN(\myifu/myicache/_1024_ ) );
AOI22_X1 \myifu/myicache/_2063_ ( .A1(\myifu/myicache/_1162_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1081_ ), .ZN(\myifu/myicache/_1025_ ) );
NAND2_X1 \myifu/myicache/_2064_ ( .A1(\myifu/myicache/_1024_ ), .A2(\myifu/myicache/_1025_ ), .ZN(\myifu/myicache/_1216_ ) );
AOI22_X1 \myifu/myicache/_2065_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1109_ ), .B1(\myifu/myicache/_0961_ ), .B2(\myifu/myicache/_1136_ ), .ZN(\myifu/myicache/_1026_ ) );
AOI22_X1 \myifu/myicache/_2066_ ( .A1(\myifu/myicache/_1163_ ), .A2(\myifu/myicache/_1003_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1082_ ), .ZN(\myifu/myicache/_1027_ ) );
NAND2_X1 \myifu/myicache/_2067_ ( .A1(\myifu/myicache/_1026_ ), .A2(\myifu/myicache/_1027_ ), .ZN(\myifu/myicache/_1217_ ) );
AOI22_X1 \myifu/myicache/_2068_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1110_ ), .B1(\myifu/myicache/_1164_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_1028_ ) );
AOI22_X1 \myifu/myicache/_2069_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1137_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1083_ ), .ZN(\myifu/myicache/_1029_ ) );
NAND2_X1 \myifu/myicache/_2070_ ( .A1(\myifu/myicache/_1028_ ), .A2(\myifu/myicache/_1029_ ), .ZN(\myifu/myicache/_1218_ ) );
AOI22_X1 \myifu/myicache/_2071_ ( .A1(\myifu/myicache/_0959_ ), .A2(\myifu/myicache/_1228_ ), .B1(\myifu/myicache/_1230_ ), .B2(\myifu/myicache/_0974_ ), .ZN(\myifu/myicache/_1030_ ) );
AOI22_X1 \myifu/myicache/_2072_ ( .A1(\myifu/myicache/_0968_ ), .A2(\myifu/myicache/_1229_ ), .B1(\myifu/myicache/_1016_ ), .B2(\myifu/myicache/_1227_ ), .ZN(\myifu/myicache/_1031_ ) );
NAND2_X1 \myifu/myicache/_2073_ ( .A1(\myifu/myicache/_1030_ ), .A2(\myifu/myicache/_1031_ ), .ZN(\myifu/myicache/_1232_ ) );
MUX2_X1 \myifu/myicache/_2074_ ( .A(\myifu/myicache/_0560_ ), .B(\myifu/myicache/_0592_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1032_ ) );
MUX2_X1 \myifu/myicache/_2075_ ( .A(\myifu/myicache/_0496_ ), .B(\myifu/myicache/_0528_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1033_ ) );
BUF_X4 \myifu/myicache/_2076_ ( .A(\myifu/myicache/_0960_ ), .Z(\myifu/myicache/_1034_ ) );
AOI22_X1 \myifu/myicache/_2077_ ( .A1(\myifu/myicache/_0974_ ), .A2(\myifu/myicache/_1032_ ), .B1(\myifu/myicache/_1033_ ), .B2(\myifu/myicache/_1034_ ), .ZN(\myifu/myicache/_1035_ ) );
INV_X1 \myifu/myicache/_2078_ ( .A(fanout_net_21 ), .ZN(\myifu/myicache/_1036_ ) );
BUF_X4 \myifu/myicache/_2079_ ( .A(\myifu/myicache/_1036_ ), .Z(\myifu/myicache/_1037_ ) );
BUF_X4 \myifu/myicache/_2080_ ( .A(\myifu/myicache/_1037_ ), .Z(\myifu/myicache/_1038_ ) );
NOR2_X1 \myifu/myicache/_2081_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0464_ ), .ZN(\myifu/myicache/_1039_ ) );
BUF_X8 \myifu/myicache/_2082_ ( .A(\myifu/myicache/_0956_ ), .Z(\myifu/myicache/_1040_ ) );
OAI211_X2 \myifu/myicache/_2083_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0432_ ), .ZN(\myifu/myicache/_1041_ ) );
NOR2_X1 \myifu/myicache/_2084_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0368_ ), .ZN(\myifu/myicache/_1042_ ) );
BUF_X4 \myifu/myicache/_2085_ ( .A(\myifu/myicache/_1037_ ), .Z(\myifu/myicache/_1043_ ) );
OAI21_X1 \myifu/myicache/_2086_ ( .A(\myifu/myicache/_1016_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0400_ ), .ZN(\myifu/myicache/_1044_ ) );
OAI221_X1 \myifu/myicache/_2087_ ( .A(\myifu/myicache/_1035_ ), .B1(\myifu/myicache/_1039_ ), .B2(\myifu/myicache/_1041_ ), .C1(\myifu/myicache/_1042_ ), .C2(\myifu/myicache/_1044_ ), .ZN(\myifu/myicache/_0656_ ) );
MUX2_X1 \myifu/myicache/_2088_ ( .A(\myifu/myicache/_0571_ ), .B(\myifu/myicache/_0603_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1045_ ) );
MUX2_X1 \myifu/myicache/_2089_ ( .A(\myifu/myicache/_0507_ ), .B(\myifu/myicache/_0539_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1046_ ) );
AOI22_X1 \myifu/myicache/_2090_ ( .A1(\myifu/myicache/_0974_ ), .A2(\myifu/myicache/_1045_ ), .B1(\myifu/myicache/_1046_ ), .B2(\myifu/myicache/_1034_ ), .ZN(\myifu/myicache/_1047_ ) );
NOR2_X1 \myifu/myicache/_2091_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0475_ ), .ZN(\myifu/myicache/_1048_ ) );
OAI211_X2 \myifu/myicache/_2092_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0443_ ), .ZN(\myifu/myicache/_1049_ ) );
NOR2_X1 \myifu/myicache/_2093_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0379_ ), .ZN(\myifu/myicache/_1050_ ) );
OAI21_X1 \myifu/myicache/_2094_ ( .A(\myifu/myicache/_1016_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0411_ ), .ZN(\myifu/myicache/_1051_ ) );
OAI221_X1 \myifu/myicache/_2095_ ( .A(\myifu/myicache/_1047_ ), .B1(\myifu/myicache/_1048_ ), .B2(\myifu/myicache/_1049_ ), .C1(\myifu/myicache/_1050_ ), .C2(\myifu/myicache/_1051_ ), .ZN(\myifu/myicache/_0667_ ) );
BUF_X4 \myifu/myicache/_2096_ ( .A(\myifu/myicache/_0971_ ), .Z(\myifu/myicache/_1052_ ) );
MUX2_X1 \myifu/myicache/_2097_ ( .A(\myifu/myicache/_0582_ ), .B(\myifu/myicache/_0614_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1053_ ) );
MUX2_X1 \myifu/myicache/_2098_ ( .A(\myifu/myicache/_0518_ ), .B(\myifu/myicache/_0550_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1054_ ) );
AOI22_X1 \myifu/myicache/_2099_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_1053_ ), .B1(\myifu/myicache/_1054_ ), .B2(\myifu/myicache/_1034_ ), .ZN(\myifu/myicache/_1055_ ) );
NOR2_X1 \myifu/myicache/_2100_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0486_ ), .ZN(\myifu/myicache/_1056_ ) );
OAI211_X2 \myifu/myicache/_2101_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0454_ ), .ZN(\myifu/myicache/_1057_ ) );
NOR2_X1 \myifu/myicache/_2102_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0390_ ), .ZN(\myifu/myicache/_1058_ ) );
BUF_X4 \myifu/myicache/_2103_ ( .A(\myifu/myicache/_0963_ ), .Z(\myifu/myicache/_1059_ ) );
OAI21_X1 \myifu/myicache/_2104_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0422_ ), .ZN(\myifu/myicache/_1060_ ) );
OAI221_X1 \myifu/myicache/_2105_ ( .A(\myifu/myicache/_1055_ ), .B1(\myifu/myicache/_1056_ ), .B2(\myifu/myicache/_1057_ ), .C1(\myifu/myicache/_1058_ ), .C2(\myifu/myicache/_1060_ ), .ZN(\myifu/myicache/_0678_ ) );
MUX2_X1 \myifu/myicache/_2106_ ( .A(\myifu/myicache/_0585_ ), .B(\myifu/myicache/_0617_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1061_ ) );
MUX2_X1 \myifu/myicache/_2107_ ( .A(\myifu/myicache/_0521_ ), .B(\myifu/myicache/_0553_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_1062_ ) );
AOI22_X1 \myifu/myicache/_2108_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_1061_ ), .B1(\myifu/myicache/_1062_ ), .B2(\myifu/myicache/_1034_ ), .ZN(\myifu/myicache/_0690_ ) );
NOR2_X1 \myifu/myicache/_2109_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0489_ ), .ZN(\myifu/myicache/_0691_ ) );
OAI211_X2 \myifu/myicache/_2110_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0457_ ), .ZN(\myifu/myicache/_0692_ ) );
NOR2_X1 \myifu/myicache/_2111_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0393_ ), .ZN(\myifu/myicache/_0693_ ) );
OAI21_X1 \myifu/myicache/_2112_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0425_ ), .ZN(\myifu/myicache/_0694_ ) );
OAI221_X1 \myifu/myicache/_2113_ ( .A(\myifu/myicache/_0690_ ), .B1(\myifu/myicache/_0691_ ), .B2(\myifu/myicache/_0692_ ), .C1(\myifu/myicache/_0693_ ), .C2(\myifu/myicache/_0694_ ), .ZN(\myifu/myicache/_0681_ ) );
MUX2_X1 \myifu/myicache/_2114_ ( .A(\myifu/myicache/_0586_ ), .B(\myifu/myicache/_0618_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0695_ ) );
MUX2_X1 \myifu/myicache/_2115_ ( .A(\myifu/myicache/_0522_ ), .B(\myifu/myicache/_0554_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0696_ ) );
AOI22_X1 \myifu/myicache/_2116_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0695_ ), .B1(\myifu/myicache/_0696_ ), .B2(\myifu/myicache/_1034_ ), .ZN(\myifu/myicache/_0697_ ) );
NOR2_X1 \myifu/myicache/_2117_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0490_ ), .ZN(\myifu/myicache/_0698_ ) );
OAI211_X2 \myifu/myicache/_2118_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0458_ ), .ZN(\myifu/myicache/_0699_ ) );
NOR2_X1 \myifu/myicache/_2119_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0394_ ), .ZN(\myifu/myicache/_0700_ ) );
OAI21_X1 \myifu/myicache/_2120_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0426_ ), .ZN(\myifu/myicache/_0701_ ) );
OAI221_X1 \myifu/myicache/_2121_ ( .A(\myifu/myicache/_0697_ ), .B1(\myifu/myicache/_0698_ ), .B2(\myifu/myicache/_0699_ ), .C1(\myifu/myicache/_0700_ ), .C2(\myifu/myicache/_0701_ ), .ZN(\myifu/myicache/_0682_ ) );
MUX2_X1 \myifu/myicache/_2122_ ( .A(\myifu/myicache/_0587_ ), .B(\myifu/myicache/_0619_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0702_ ) );
MUX2_X1 \myifu/myicache/_2123_ ( .A(\myifu/myicache/_0459_ ), .B(\myifu/myicache/_0491_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0703_ ) );
AOI22_X1 \myifu/myicache/_2124_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0702_ ), .B1(\myifu/myicache/_0703_ ), .B2(\myifu/myicache/_0959_ ), .ZN(\myifu/myicache/_0704_ ) );
NOR2_X1 \myifu/myicache/_2125_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0523_ ), .ZN(\myifu/myicache/_0705_ ) );
OAI21_X1 \myifu/myicache/_2126_ ( .A(\myifu/myicache/_1034_ ), .B1(\myifu/myicache/_1037_ ), .B2(\myifu/myicache/_0555_ ), .ZN(\myifu/myicache/_0706_ ) );
NOR2_X1 \myifu/myicache/_2127_ ( .A1(fanout_net_21 ), .A2(\myifu/myicache/_0395_ ), .ZN(\myifu/myicache/_0707_ ) );
OAI21_X1 \myifu/myicache/_2128_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0427_ ), .ZN(\myifu/myicache/_0708_ ) );
OAI221_X1 \myifu/myicache/_2129_ ( .A(\myifu/myicache/_0704_ ), .B1(\myifu/myicache/_0705_ ), .B2(\myifu/myicache/_0706_ ), .C1(\myifu/myicache/_0707_ ), .C2(\myifu/myicache/_0708_ ), .ZN(\myifu/myicache/_0683_ ) );
BUF_X4 \myifu/myicache/_2130_ ( .A(\myifu/myicache/_0963_ ), .Z(\myifu/myicache/_0709_ ) );
MUX2_X1 \myifu/myicache/_2131_ ( .A(\myifu/myicache/_0396_ ), .B(\myifu/myicache/_0428_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0710_ ) );
MUX2_X1 \myifu/myicache/_2132_ ( .A(\myifu/myicache/_0524_ ), .B(\myifu/myicache/_0556_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0711_ ) );
BUF_X4 \myifu/myicache/_2133_ ( .A(\myifu/myicache/_0960_ ), .Z(\myifu/myicache/_0712_ ) );
AOI22_X1 \myifu/myicache/_2134_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0710_ ), .B1(\myifu/myicache/_0711_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0713_ ) );
NOR2_X1 \myifu/myicache/_2135_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0620_ ), .ZN(\myifu/myicache/_0714_ ) );
OAI211_X2 \myifu/myicache/_2136_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0588_ ), .ZN(\myifu/myicache/_0715_ ) );
BUF_X4 \myifu/myicache/_2137_ ( .A(\myifu/myicache/_1037_ ), .Z(\myifu/myicache/_0716_ ) );
NOR2_X1 \myifu/myicache/_2138_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0492_ ), .ZN(\myifu/myicache/_0717_ ) );
BUF_X8 \myifu/myicache/_2139_ ( .A(\myifu/myicache/_0956_ ), .Z(\myifu/myicache/_0718_ ) );
OAI211_X2 \myifu/myicache/_2140_ ( .A(\myifu/myicache/_0718_ ), .B(fanout_net_20 ), .C1(fanout_net_21 ), .C2(\myifu/myicache/_0460_ ), .ZN(\myifu/myicache/_0719_ ) );
OAI221_X1 \myifu/myicache/_2141_ ( .A(\myifu/myicache/_0713_ ), .B1(\myifu/myicache/_0714_ ), .B2(\myifu/myicache/_0715_ ), .C1(\myifu/myicache/_0717_ ), .C2(\myifu/myicache/_0719_ ), .ZN(\myifu/myicache/_0684_ ) );
MUX2_X1 \myifu/myicache/_2142_ ( .A(\myifu/myicache/_0589_ ), .B(\myifu/myicache/_0621_ ), .S(fanout_net_21 ), .Z(\myifu/myicache/_0720_ ) );
MUX2_X1 \myifu/myicache/_2143_ ( .A(\myifu/myicache/_0525_ ), .B(\myifu/myicache/_0557_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0721_ ) );
AOI22_X1 \myifu/myicache/_2144_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0720_ ), .B1(\myifu/myicache/_0721_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0722_ ) );
NOR2_X1 \myifu/myicache/_2145_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0493_ ), .ZN(\myifu/myicache/_0723_ ) );
OAI211_X2 \myifu/myicache/_2146_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0461_ ), .ZN(\myifu/myicache/_0724_ ) );
NOR2_X1 \myifu/myicache/_2147_ ( .A1(fanout_net_22 ), .A2(\myifu/myicache/_0397_ ), .ZN(\myifu/myicache/_0725_ ) );
OAI21_X1 \myifu/myicache/_2148_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0429_ ), .ZN(\myifu/myicache/_0726_ ) );
OAI221_X1 \myifu/myicache/_2149_ ( .A(\myifu/myicache/_0722_ ), .B1(\myifu/myicache/_0723_ ), .B2(\myifu/myicache/_0724_ ), .C1(\myifu/myicache/_0725_ ), .C2(\myifu/myicache/_0726_ ), .ZN(\myifu/myicache/_0685_ ) );
MUX2_X1 \myifu/myicache/_2150_ ( .A(\myifu/myicache/_0590_ ), .B(\myifu/myicache/_0622_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0727_ ) );
MUX2_X1 \myifu/myicache/_2151_ ( .A(\myifu/myicache/_0526_ ), .B(\myifu/myicache/_0558_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0728_ ) );
AOI22_X1 \myifu/myicache/_2152_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0727_ ), .B1(\myifu/myicache/_0728_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0729_ ) );
NOR2_X1 \myifu/myicache/_2153_ ( .A1(\myifu/myicache/_1038_ ), .A2(\myifu/myicache/_0494_ ), .ZN(\myifu/myicache/_0730_ ) );
OAI211_X2 \myifu/myicache/_2154_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0462_ ), .ZN(\myifu/myicache/_0731_ ) );
NOR2_X1 \myifu/myicache/_2155_ ( .A1(fanout_net_22 ), .A2(\myifu/myicache/_0398_ ), .ZN(\myifu/myicache/_0732_ ) );
OAI21_X1 \myifu/myicache/_2156_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_1043_ ), .B2(\myifu/myicache/_0430_ ), .ZN(\myifu/myicache/_0733_ ) );
OAI221_X1 \myifu/myicache/_2157_ ( .A(\myifu/myicache/_0729_ ), .B1(\myifu/myicache/_0730_ ), .B2(\myifu/myicache/_0731_ ), .C1(\myifu/myicache/_0732_ ), .C2(\myifu/myicache/_0733_ ), .ZN(\myifu/myicache/_0686_ ) );
MUX2_X1 \myifu/myicache/_2158_ ( .A(\myifu/myicache/_0591_ ), .B(\myifu/myicache/_0623_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0734_ ) );
MUX2_X1 \myifu/myicache/_2159_ ( .A(\myifu/myicache/_0527_ ), .B(\myifu/myicache/_0559_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0735_ ) );
AOI22_X1 \myifu/myicache/_2160_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0734_ ), .B1(\myifu/myicache/_0735_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0736_ ) );
BUF_X4 \myifu/myicache/_2161_ ( .A(\myifu/myicache/_1037_ ), .Z(\myifu/myicache/_0737_ ) );
NOR2_X1 \myifu/myicache/_2162_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0495_ ), .ZN(\myifu/myicache/_0738_ ) );
OAI211_X2 \myifu/myicache/_2163_ ( .A(\myifu/myicache/_1040_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0463_ ), .ZN(\myifu/myicache/_0739_ ) );
NOR2_X1 \myifu/myicache/_2164_ ( .A1(fanout_net_22 ), .A2(\myifu/myicache/_0399_ ), .ZN(\myifu/myicache/_0740_ ) );
BUF_X4 \myifu/myicache/_2165_ ( .A(\myifu/myicache/_1037_ ), .Z(\myifu/myicache/_0741_ ) );
OAI21_X1 \myifu/myicache/_2166_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0431_ ), .ZN(\myifu/myicache/_0742_ ) );
OAI221_X1 \myifu/myicache/_2167_ ( .A(\myifu/myicache/_0736_ ), .B1(\myifu/myicache/_0738_ ), .B2(\myifu/myicache/_0739_ ), .C1(\myifu/myicache/_0740_ ), .C2(\myifu/myicache/_0742_ ), .ZN(\myifu/myicache/_0687_ ) );
MUX2_X1 \myifu/myicache/_2168_ ( .A(\myifu/myicache/_0369_ ), .B(\myifu/myicache/_0401_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0743_ ) );
MUX2_X1 \myifu/myicache/_2169_ ( .A(\myifu/myicache/_0497_ ), .B(\myifu/myicache/_0529_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0744_ ) );
AOI22_X1 \myifu/myicache/_2170_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0743_ ), .B1(\myifu/myicache/_0744_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0745_ ) );
NOR2_X1 \myifu/myicache/_2171_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0593_ ), .ZN(\myifu/myicache/_0746_ ) );
OAI211_X2 \myifu/myicache/_2172_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0561_ ), .ZN(\myifu/myicache/_0747_ ) );
NOR2_X1 \myifu/myicache/_2173_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0465_ ), .ZN(\myifu/myicache/_0748_ ) );
OAI211_X2 \myifu/myicache/_2174_ ( .A(\myifu/myicache/_0718_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0433_ ), .ZN(\myifu/myicache/_0749_ ) );
OAI221_X1 \myifu/myicache/_2175_ ( .A(\myifu/myicache/_0745_ ), .B1(\myifu/myicache/_0746_ ), .B2(\myifu/myicache/_0747_ ), .C1(\myifu/myicache/_0748_ ), .C2(\myifu/myicache/_0749_ ), .ZN(\myifu/myicache/_0657_ ) );
MUX2_X1 \myifu/myicache/_2176_ ( .A(\myifu/myicache/_0562_ ), .B(\myifu/myicache/_0594_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0750_ ) );
MUX2_X1 \myifu/myicache/_2177_ ( .A(\myifu/myicache/_0498_ ), .B(\myifu/myicache/_0530_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0751_ ) );
AOI22_X1 \myifu/myicache/_2178_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0750_ ), .B1(\myifu/myicache/_0751_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0752_ ) );
NOR2_X1 \myifu/myicache/_2179_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0466_ ), .ZN(\myifu/myicache/_0753_ ) );
OAI211_X2 \myifu/myicache/_2180_ ( .A(\myifu/myicache/_0956_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0434_ ), .ZN(\myifu/myicache/_0754_ ) );
NOR2_X1 \myifu/myicache/_2181_ ( .A1(fanout_net_22 ), .A2(\myifu/myicache/_0370_ ), .ZN(\myifu/myicache/_0755_ ) );
OAI21_X1 \myifu/myicache/_2182_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0402_ ), .ZN(\myifu/myicache/_0756_ ) );
OAI221_X1 \myifu/myicache/_2183_ ( .A(\myifu/myicache/_0752_ ), .B1(\myifu/myicache/_0753_ ), .B2(\myifu/myicache/_0754_ ), .C1(\myifu/myicache/_0755_ ), .C2(\myifu/myicache/_0756_ ), .ZN(\myifu/myicache/_0658_ ) );
MUX2_X1 \myifu/myicache/_2184_ ( .A(\myifu/myicache/_0371_ ), .B(\myifu/myicache/_0403_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0757_ ) );
MUX2_X1 \myifu/myicache/_2185_ ( .A(\myifu/myicache/_0435_ ), .B(\myifu/myicache/_0467_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0758_ ) );
AOI22_X1 \myifu/myicache/_2186_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0757_ ), .B1(\myifu/myicache/_0758_ ), .B2(\myifu/myicache/_0959_ ), .ZN(\myifu/myicache/_0759_ ) );
NOR2_X1 \myifu/myicache/_2187_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0595_ ), .ZN(\myifu/myicache/_0760_ ) );
OAI211_X2 \myifu/myicache/_2188_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0563_ ), .ZN(\myifu/myicache/_0761_ ) );
NOR2_X1 \myifu/myicache/_2189_ ( .A1(fanout_net_22 ), .A2(\myifu/myicache/_0499_ ), .ZN(\myifu/myicache/_0762_ ) );
OAI21_X1 \myifu/myicache/_2190_ ( .A(\myifu/myicache/_0961_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0531_ ), .ZN(\myifu/myicache/_0763_ ) );
OAI221_X1 \myifu/myicache/_2191_ ( .A(\myifu/myicache/_0759_ ), .B1(\myifu/myicache/_0760_ ), .B2(\myifu/myicache/_0761_ ), .C1(\myifu/myicache/_0762_ ), .C2(\myifu/myicache/_0763_ ), .ZN(\myifu/myicache/_0659_ ) );
MUX2_X1 \myifu/myicache/_2192_ ( .A(\myifu/myicache/_0372_ ), .B(\myifu/myicache/_0404_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0764_ ) );
MUX2_X1 \myifu/myicache/_2193_ ( .A(\myifu/myicache/_0500_ ), .B(\myifu/myicache/_0532_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0765_ ) );
AOI22_X1 \myifu/myicache/_2194_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0764_ ), .B1(\myifu/myicache/_0765_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0766_ ) );
NOR2_X1 \myifu/myicache/_2195_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0596_ ), .ZN(\myifu/myicache/_0767_ ) );
OAI211_X2 \myifu/myicache/_2196_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0564_ ), .ZN(\myifu/myicache/_0768_ ) );
NOR2_X1 \myifu/myicache/_2197_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0468_ ), .ZN(\myifu/myicache/_0769_ ) );
OAI211_X2 \myifu/myicache/_2198_ ( .A(\myifu/myicache/_0718_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0436_ ), .ZN(\myifu/myicache/_0770_ ) );
OAI221_X1 \myifu/myicache/_2199_ ( .A(\myifu/myicache/_0766_ ), .B1(\myifu/myicache/_0767_ ), .B2(\myifu/myicache/_0768_ ), .C1(\myifu/myicache/_0769_ ), .C2(\myifu/myicache/_0770_ ), .ZN(\myifu/myicache/_0660_ ) );
MUX2_X1 \myifu/myicache/_2200_ ( .A(\myifu/myicache/_0565_ ), .B(\myifu/myicache/_0597_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0771_ ) );
MUX2_X1 \myifu/myicache/_2201_ ( .A(\myifu/myicache/_0501_ ), .B(\myifu/myicache/_0533_ ), .S(fanout_net_22 ), .Z(\myifu/myicache/_0772_ ) );
AOI22_X1 \myifu/myicache/_2202_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0771_ ), .B1(\myifu/myicache/_0772_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0773_ ) );
NOR2_X1 \myifu/myicache/_2203_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0469_ ), .ZN(\myifu/myicache/_0774_ ) );
OAI211_X2 \myifu/myicache/_2204_ ( .A(\myifu/myicache/_0956_ ), .B(fanout_net_20 ), .C1(fanout_net_22 ), .C2(\myifu/myicache/_0437_ ), .ZN(\myifu/myicache/_0775_ ) );
NOR2_X1 \myifu/myicache/_2205_ ( .A1(fanout_net_23 ), .A2(\myifu/myicache/_0373_ ), .ZN(\myifu/myicache/_0776_ ) );
OAI21_X1 \myifu/myicache/_2206_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0405_ ), .ZN(\myifu/myicache/_0777_ ) );
OAI221_X1 \myifu/myicache/_2207_ ( .A(\myifu/myicache/_0773_ ), .B1(\myifu/myicache/_0774_ ), .B2(\myifu/myicache/_0775_ ), .C1(\myifu/myicache/_0776_ ), .C2(\myifu/myicache/_0777_ ), .ZN(\myifu/myicache/_0661_ ) );
MUX2_X1 \myifu/myicache/_2208_ ( .A(\myifu/myicache/_0374_ ), .B(\myifu/myicache/_0406_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0778_ ) );
MUX2_X1 \myifu/myicache/_2209_ ( .A(\myifu/myicache/_0502_ ), .B(\myifu/myicache/_0534_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0779_ ) );
AOI22_X1 \myifu/myicache/_2210_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0778_ ), .B1(\myifu/myicache/_0779_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0780_ ) );
NOR2_X1 \myifu/myicache/_2211_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0598_ ), .ZN(\myifu/myicache/_0781_ ) );
OAI211_X2 \myifu/myicache/_2212_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0566_ ), .ZN(\myifu/myicache/_0782_ ) );
NOR2_X1 \myifu/myicache/_2213_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0470_ ), .ZN(\myifu/myicache/_0783_ ) );
OAI211_X2 \myifu/myicache/_2214_ ( .A(\myifu/myicache/_0718_ ), .B(fanout_net_20 ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0438_ ), .ZN(\myifu/myicache/_0784_ ) );
OAI221_X1 \myifu/myicache/_2215_ ( .A(\myifu/myicache/_0780_ ), .B1(\myifu/myicache/_0781_ ), .B2(\myifu/myicache/_0782_ ), .C1(\myifu/myicache/_0783_ ), .C2(\myifu/myicache/_0784_ ), .ZN(\myifu/myicache/_0662_ ) );
MUX2_X1 \myifu/myicache/_2216_ ( .A(\myifu/myicache/_0375_ ), .B(\myifu/myicache/_0407_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0785_ ) );
MUX2_X1 \myifu/myicache/_2217_ ( .A(\myifu/myicache/_0503_ ), .B(\myifu/myicache/_0535_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0786_ ) );
AOI22_X1 \myifu/myicache/_2218_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0785_ ), .B1(\myifu/myicache/_0786_ ), .B2(\myifu/myicache/_0712_ ), .ZN(\myifu/myicache/_0787_ ) );
NOR2_X1 \myifu/myicache/_2219_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0599_ ), .ZN(\myifu/myicache/_0788_ ) );
OAI211_X2 \myifu/myicache/_2220_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0567_ ), .ZN(\myifu/myicache/_0789_ ) );
NOR2_X1 \myifu/myicache/_2221_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0471_ ), .ZN(\myifu/myicache/_0790_ ) );
OAI211_X2 \myifu/myicache/_2222_ ( .A(\myifu/myicache/_0718_ ), .B(fanout_net_20 ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0439_ ), .ZN(\myifu/myicache/_0791_ ) );
OAI221_X1 \myifu/myicache/_2223_ ( .A(\myifu/myicache/_0787_ ), .B1(\myifu/myicache/_0788_ ), .B2(\myifu/myicache/_0789_ ), .C1(\myifu/myicache/_0790_ ), .C2(\myifu/myicache/_0791_ ), .ZN(\myifu/myicache/_0663_ ) );
MUX2_X1 \myifu/myicache/_2224_ ( .A(\myifu/myicache/_0568_ ), .B(\myifu/myicache/_0600_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0792_ ) );
MUX2_X1 \myifu/myicache/_2225_ ( .A(\myifu/myicache/_0504_ ), .B(\myifu/myicache/_0536_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0793_ ) );
BUF_X4 \myifu/myicache/_2226_ ( .A(\myifu/myicache/_0960_ ), .Z(\myifu/myicache/_0794_ ) );
AOI22_X1 \myifu/myicache/_2227_ ( .A1(\myifu/myicache/_1052_ ), .A2(\myifu/myicache/_0792_ ), .B1(\myifu/myicache/_0793_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0795_ ) );
NOR2_X1 \myifu/myicache/_2228_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0472_ ), .ZN(\myifu/myicache/_0796_ ) );
OAI211_X2 \myifu/myicache/_2229_ ( .A(\myifu/myicache/_0956_ ), .B(fanout_net_20 ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0440_ ), .ZN(\myifu/myicache/_0797_ ) );
NOR2_X1 \myifu/myicache/_2230_ ( .A1(fanout_net_23 ), .A2(\myifu/myicache/_0376_ ), .ZN(\myifu/myicache/_0798_ ) );
OAI21_X1 \myifu/myicache/_2231_ ( .A(\myifu/myicache/_1059_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0408_ ), .ZN(\myifu/myicache/_0799_ ) );
OAI221_X1 \myifu/myicache/_2232_ ( .A(\myifu/myicache/_0795_ ), .B1(\myifu/myicache/_0796_ ), .B2(\myifu/myicache/_0797_ ), .C1(\myifu/myicache/_0798_ ), .C2(\myifu/myicache/_0799_ ), .ZN(\myifu/myicache/_0664_ ) );
MUX2_X1 \myifu/myicache/_2233_ ( .A(\myifu/myicache/_0569_ ), .B(\myifu/myicache/_0601_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0800_ ) );
MUX2_X1 \myifu/myicache/_2234_ ( .A(\myifu/myicache/_0505_ ), .B(\myifu/myicache/_0537_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0801_ ) );
AOI22_X1 \myifu/myicache/_2235_ ( .A1(\myifu/myicache/_0971_ ), .A2(\myifu/myicache/_0800_ ), .B1(\myifu/myicache/_0801_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0802_ ) );
NOR2_X1 \myifu/myicache/_2236_ ( .A1(\myifu/myicache/_0737_ ), .A2(\myifu/myicache/_0473_ ), .ZN(\myifu/myicache/_0803_ ) );
OAI211_X2 \myifu/myicache/_2237_ ( .A(\myifu/myicache/_0956_ ), .B(fanout_net_20 ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0441_ ), .ZN(\myifu/myicache/_0804_ ) );
NOR2_X1 \myifu/myicache/_2238_ ( .A1(fanout_net_23 ), .A2(\myifu/myicache/_0377_ ), .ZN(\myifu/myicache/_0805_ ) );
OAI21_X1 \myifu/myicache/_2239_ ( .A(\myifu/myicache/_0709_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0409_ ), .ZN(\myifu/myicache/_0806_ ) );
OAI221_X1 \myifu/myicache/_2240_ ( .A(\myifu/myicache/_0802_ ), .B1(\myifu/myicache/_0803_ ), .B2(\myifu/myicache/_0804_ ), .C1(\myifu/myicache/_0805_ ), .C2(\myifu/myicache/_0806_ ), .ZN(\myifu/myicache/_0665_ ) );
MUX2_X1 \myifu/myicache/_2241_ ( .A(\myifu/myicache/_0378_ ), .B(\myifu/myicache/_0410_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0807_ ) );
MUX2_X1 \myifu/myicache/_2242_ ( .A(\myifu/myicache/_0506_ ), .B(\myifu/myicache/_0538_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0808_ ) );
AOI22_X1 \myifu/myicache/_2243_ ( .A1(\myifu/myicache/_0709_ ), .A2(\myifu/myicache/_0807_ ), .B1(\myifu/myicache/_0808_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0809_ ) );
BUF_X4 \myifu/myicache/_2244_ ( .A(\myifu/myicache/_1037_ ), .Z(\myifu/myicache/_0810_ ) );
NOR2_X1 \myifu/myicache/_2245_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0602_ ), .ZN(\myifu/myicache/_0811_ ) );
OAI211_X2 \myifu/myicache/_2246_ ( .A(fanout_net_20 ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0570_ ), .ZN(\myifu/myicache/_0812_ ) );
NOR2_X1 \myifu/myicache/_2247_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0474_ ), .ZN(\myifu/myicache/_0813_ ) );
OAI211_X2 \myifu/myicache/_2248_ ( .A(\myifu/myicache/_0718_ ), .B(fanout_net_20 ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0442_ ), .ZN(\myifu/myicache/_0814_ ) );
OAI221_X1 \myifu/myicache/_2249_ ( .A(\myifu/myicache/_0809_ ), .B1(\myifu/myicache/_0811_ ), .B2(\myifu/myicache/_0812_ ), .C1(\myifu/myicache/_0813_ ), .C2(\myifu/myicache/_0814_ ), .ZN(\myifu/myicache/_0666_ ) );
BUF_X4 \myifu/myicache/_2250_ ( .A(\myifu/myicache/_0963_ ), .Z(\myifu/myicache/_0815_ ) );
MUX2_X1 \myifu/myicache/_2251_ ( .A(\myifu/myicache/_0380_ ), .B(\myifu/myicache/_0412_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0816_ ) );
MUX2_X1 \myifu/myicache/_2252_ ( .A(\myifu/myicache/_0444_ ), .B(\myifu/myicache/_0476_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0817_ ) );
AOI22_X1 \myifu/myicache/_2253_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0816_ ), .B1(\myifu/myicache/_0817_ ), .B2(\myifu/myicache/_0958_ ), .ZN(\myifu/myicache/_0818_ ) );
NOR2_X1 \myifu/myicache/_2254_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0604_ ), .ZN(\myifu/myicache/_0819_ ) );
OAI211_X2 \myifu/myicache/_2255_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_23 ), .C2(\myifu/myicache/_0572_ ), .ZN(\myifu/myicache/_0820_ ) );
NOR2_X1 \myifu/myicache/_2256_ ( .A1(fanout_net_23 ), .A2(\myifu/myicache/_0508_ ), .ZN(\myifu/myicache/_0821_ ) );
OAI21_X1 \myifu/myicache/_2257_ ( .A(\myifu/myicache/_0961_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0540_ ), .ZN(\myifu/myicache/_0822_ ) );
OAI221_X1 \myifu/myicache/_2258_ ( .A(\myifu/myicache/_0818_ ), .B1(\myifu/myicache/_0819_ ), .B2(\myifu/myicache/_0820_ ), .C1(\myifu/myicache/_0821_ ), .C2(\myifu/myicache/_0822_ ), .ZN(\myifu/myicache/_0668_ ) );
MUX2_X1 \myifu/myicache/_2259_ ( .A(\myifu/myicache/_0573_ ), .B(\myifu/myicache/_0605_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0823_ ) );
MUX2_X1 \myifu/myicache/_2260_ ( .A(\myifu/myicache/_0445_ ), .B(\myifu/myicache/_0477_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0824_ ) );
AOI22_X1 \myifu/myicache/_2261_ ( .A1(\myifu/myicache/_0971_ ), .A2(\myifu/myicache/_0823_ ), .B1(\myifu/myicache/_0824_ ), .B2(\myifu/myicache/_0958_ ), .ZN(\myifu/myicache/_0825_ ) );
NOR2_X1 \myifu/myicache/_2262_ ( .A1(fanout_net_23 ), .A2(\myifu/myicache/_0509_ ), .ZN(\myifu/myicache/_0826_ ) );
OAI21_X1 \myifu/myicache/_2263_ ( .A(\myifu/myicache/_1034_ ), .B1(\myifu/myicache/_1037_ ), .B2(\myifu/myicache/_0541_ ), .ZN(\myifu/myicache/_0827_ ) );
NOR2_X1 \myifu/myicache/_2264_ ( .A1(fanout_net_23 ), .A2(\myifu/myicache/_0381_ ), .ZN(\myifu/myicache/_0828_ ) );
OAI21_X1 \myifu/myicache/_2265_ ( .A(\myifu/myicache/_0709_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0413_ ), .ZN(\myifu/myicache/_0829_ ) );
OAI221_X1 \myifu/myicache/_2266_ ( .A(\myifu/myicache/_0825_ ), .B1(\myifu/myicache/_0826_ ), .B2(\myifu/myicache/_0827_ ), .C1(\myifu/myicache/_0828_ ), .C2(\myifu/myicache/_0829_ ), .ZN(\myifu/myicache/_0669_ ) );
MUX2_X1 \myifu/myicache/_2267_ ( .A(\myifu/myicache/_0382_ ), .B(\myifu/myicache/_0414_ ), .S(fanout_net_23 ), .Z(\myifu/myicache/_0830_ ) );
MUX2_X1 \myifu/myicache/_2268_ ( .A(\myifu/myicache/_0510_ ), .B(\myifu/myicache/_0542_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0831_ ) );
AOI22_X1 \myifu/myicache/_2269_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0830_ ), .B1(\myifu/myicache/_0831_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0832_ ) );
NOR2_X1 \myifu/myicache/_2270_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0606_ ), .ZN(\myifu/myicache/_0833_ ) );
OAI211_X2 \myifu/myicache/_2271_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0574_ ), .ZN(\myifu/myicache/_0834_ ) );
NOR2_X1 \myifu/myicache/_2272_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0478_ ), .ZN(\myifu/myicache/_0835_ ) );
OAI211_X2 \myifu/myicache/_2273_ ( .A(\myifu/myicache/_0718_ ), .B(\myifu/myicache/_0688_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0446_ ), .ZN(\myifu/myicache/_0836_ ) );
OAI221_X1 \myifu/myicache/_2274_ ( .A(\myifu/myicache/_0832_ ), .B1(\myifu/myicache/_0833_ ), .B2(\myifu/myicache/_0834_ ), .C1(\myifu/myicache/_0835_ ), .C2(\myifu/myicache/_0836_ ), .ZN(\myifu/myicache/_0670_ ) );
MUX2_X1 \myifu/myicache/_2275_ ( .A(\myifu/myicache/_0383_ ), .B(\myifu/myicache/_0415_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0837_ ) );
MUX2_X1 \myifu/myicache/_2276_ ( .A(\myifu/myicache/_0447_ ), .B(\myifu/myicache/_0479_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0838_ ) );
AOI22_X1 \myifu/myicache/_2277_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0837_ ), .B1(\myifu/myicache/_0838_ ), .B2(\myifu/myicache/_0958_ ), .ZN(\myifu/myicache/_0839_ ) );
NOR2_X1 \myifu/myicache/_2278_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0607_ ), .ZN(\myifu/myicache/_0840_ ) );
OAI211_X2 \myifu/myicache/_2279_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0575_ ), .ZN(\myifu/myicache/_0841_ ) );
NOR2_X1 \myifu/myicache/_2280_ ( .A1(fanout_net_24 ), .A2(\myifu/myicache/_0511_ ), .ZN(\myifu/myicache/_0842_ ) );
OAI21_X1 \myifu/myicache/_2281_ ( .A(\myifu/myicache/_1034_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0543_ ), .ZN(\myifu/myicache/_0843_ ) );
OAI221_X1 \myifu/myicache/_2282_ ( .A(\myifu/myicache/_0839_ ), .B1(\myifu/myicache/_0840_ ), .B2(\myifu/myicache/_0841_ ), .C1(\myifu/myicache/_0842_ ), .C2(\myifu/myicache/_0843_ ), .ZN(\myifu/myicache/_0671_ ) );
MUX2_X1 \myifu/myicache/_2283_ ( .A(\myifu/myicache/_0384_ ), .B(\myifu/myicache/_0416_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0844_ ) );
MUX2_X1 \myifu/myicache/_2284_ ( .A(\myifu/myicache/_0512_ ), .B(\myifu/myicache/_0544_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0845_ ) );
AOI22_X1 \myifu/myicache/_2285_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0844_ ), .B1(\myifu/myicache/_0845_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0846_ ) );
NOR2_X1 \myifu/myicache/_2286_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0608_ ), .ZN(\myifu/myicache/_0847_ ) );
OAI211_X2 \myifu/myicache/_2287_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0576_ ), .ZN(\myifu/myicache/_0848_ ) );
NOR2_X1 \myifu/myicache/_2288_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0480_ ), .ZN(\myifu/myicache/_0849_ ) );
OAI211_X2 \myifu/myicache/_2289_ ( .A(\myifu/myicache/_0718_ ), .B(\myifu/myicache/_0688_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0448_ ), .ZN(\myifu/myicache/_0850_ ) );
OAI221_X1 \myifu/myicache/_2290_ ( .A(\myifu/myicache/_0846_ ), .B1(\myifu/myicache/_0847_ ), .B2(\myifu/myicache/_0848_ ), .C1(\myifu/myicache/_0849_ ), .C2(\myifu/myicache/_0850_ ), .ZN(\myifu/myicache/_0672_ ) );
MUX2_X1 \myifu/myicache/_2291_ ( .A(\myifu/myicache/_0385_ ), .B(\myifu/myicache/_0417_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0851_ ) );
MUX2_X1 \myifu/myicache/_2292_ ( .A(\myifu/myicache/_0513_ ), .B(\myifu/myicache/_0545_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0852_ ) );
AOI22_X1 \myifu/myicache/_2293_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0851_ ), .B1(\myifu/myicache/_0852_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0853_ ) );
NOR2_X1 \myifu/myicache/_2294_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0609_ ), .ZN(\myifu/myicache/_0854_ ) );
OAI211_X2 \myifu/myicache/_2295_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0577_ ), .ZN(\myifu/myicache/_0855_ ) );
NOR2_X1 \myifu/myicache/_2296_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0481_ ), .ZN(\myifu/myicache/_0856_ ) );
OAI211_X2 \myifu/myicache/_2297_ ( .A(\myifu/myicache/_0718_ ), .B(\myifu/myicache/_0688_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0449_ ), .ZN(\myifu/myicache/_0857_ ) );
OAI221_X1 \myifu/myicache/_2298_ ( .A(\myifu/myicache/_0853_ ), .B1(\myifu/myicache/_0854_ ), .B2(\myifu/myicache/_0855_ ), .C1(\myifu/myicache/_0856_ ), .C2(\myifu/myicache/_0857_ ), .ZN(\myifu/myicache/_0673_ ) );
MUX2_X1 \myifu/myicache/_2299_ ( .A(\myifu/myicache/_0386_ ), .B(\myifu/myicache/_0418_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0858_ ) );
MUX2_X1 \myifu/myicache/_2300_ ( .A(\myifu/myicache/_0450_ ), .B(\myifu/myicache/_0482_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0859_ ) );
AOI22_X1 \myifu/myicache/_2301_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0858_ ), .B1(\myifu/myicache/_0859_ ), .B2(\myifu/myicache/_0958_ ), .ZN(\myifu/myicache/_0860_ ) );
NOR2_X1 \myifu/myicache/_2302_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0610_ ), .ZN(\myifu/myicache/_0861_ ) );
OAI211_X2 \myifu/myicache/_2303_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0578_ ), .ZN(\myifu/myicache/_0862_ ) );
NOR2_X1 \myifu/myicache/_2304_ ( .A1(fanout_net_24 ), .A2(\myifu/myicache/_0514_ ), .ZN(\myifu/myicache/_0863_ ) );
OAI21_X1 \myifu/myicache/_2305_ ( .A(\myifu/myicache/_1034_ ), .B1(\myifu/myicache/_0741_ ), .B2(\myifu/myicache/_0546_ ), .ZN(\myifu/myicache/_0864_ ) );
OAI221_X1 \myifu/myicache/_2306_ ( .A(\myifu/myicache/_0860_ ), .B1(\myifu/myicache/_0861_ ), .B2(\myifu/myicache/_0862_ ), .C1(\myifu/myicache/_0863_ ), .C2(\myifu/myicache/_0864_ ), .ZN(\myifu/myicache/_0674_ ) );
MUX2_X1 \myifu/myicache/_2307_ ( .A(\myifu/myicache/_0579_ ), .B(\myifu/myicache/_0611_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0865_ ) );
MUX2_X1 \myifu/myicache/_2308_ ( .A(\myifu/myicache/_0515_ ), .B(\myifu/myicache/_0547_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0866_ ) );
AOI22_X1 \myifu/myicache/_2309_ ( .A1(\myifu/myicache/_0971_ ), .A2(\myifu/myicache/_0865_ ), .B1(\myifu/myicache/_0866_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0867_ ) );
NOR2_X1 \myifu/myicache/_2310_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0483_ ), .ZN(\myifu/myicache/_0868_ ) );
OAI211_X2 \myifu/myicache/_2311_ ( .A(\myifu/myicache/_0956_ ), .B(\myifu/myicache/_0688_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0451_ ), .ZN(\myifu/myicache/_0869_ ) );
NOR2_X1 \myifu/myicache/_2312_ ( .A1(fanout_net_24 ), .A2(\myifu/myicache/_0387_ ), .ZN(\myifu/myicache/_0870_ ) );
OAI21_X1 \myifu/myicache/_2313_ ( .A(\myifu/myicache/_0709_ ), .B1(\myifu/myicache/_1038_ ), .B2(\myifu/myicache/_0419_ ), .ZN(\myifu/myicache/_0871_ ) );
OAI221_X1 \myifu/myicache/_2314_ ( .A(\myifu/myicache/_0867_ ), .B1(\myifu/myicache/_0868_ ), .B2(\myifu/myicache/_0869_ ), .C1(\myifu/myicache/_0870_ ), .C2(\myifu/myicache/_0871_ ), .ZN(\myifu/myicache/_0675_ ) );
MUX2_X1 \myifu/myicache/_2315_ ( .A(\myifu/myicache/_0388_ ), .B(\myifu/myicache/_0420_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0872_ ) );
MUX2_X1 \myifu/myicache/_2316_ ( .A(\myifu/myicache/_0516_ ), .B(\myifu/myicache/_0548_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0873_ ) );
AOI22_X1 \myifu/myicache/_2317_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0872_ ), .B1(\myifu/myicache/_0873_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0874_ ) );
NOR2_X1 \myifu/myicache/_2318_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0612_ ), .ZN(\myifu/myicache/_0875_ ) );
OAI211_X2 \myifu/myicache/_2319_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0580_ ), .ZN(\myifu/myicache/_0876_ ) );
NOR2_X1 \myifu/myicache/_2320_ ( .A1(\myifu/myicache/_0716_ ), .A2(\myifu/myicache/_0484_ ), .ZN(\myifu/myicache/_0877_ ) );
OAI211_X2 \myifu/myicache/_2321_ ( .A(\myifu/myicache/_0718_ ), .B(\myifu/myicache/_0688_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0452_ ), .ZN(\myifu/myicache/_0878_ ) );
OAI221_X1 \myifu/myicache/_2322_ ( .A(\myifu/myicache/_0874_ ), .B1(\myifu/myicache/_0875_ ), .B2(\myifu/myicache/_0876_ ), .C1(\myifu/myicache/_0877_ ), .C2(\myifu/myicache/_0878_ ), .ZN(\myifu/myicache/_0676_ ) );
MUX2_X1 \myifu/myicache/_2323_ ( .A(\myifu/myicache/_0389_ ), .B(\myifu/myicache/_0421_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0879_ ) );
MUX2_X1 \myifu/myicache/_2324_ ( .A(\myifu/myicache/_0453_ ), .B(\myifu/myicache/_0485_ ), .S(fanout_net_24 ), .Z(\myifu/myicache/_0880_ ) );
AOI22_X1 \myifu/myicache/_2325_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0879_ ), .B1(\myifu/myicache/_0880_ ), .B2(\myifu/myicache/_0958_ ), .ZN(\myifu/myicache/_0881_ ) );
NOR2_X1 \myifu/myicache/_2326_ ( .A1(\myifu/myicache/_0810_ ), .A2(\myifu/myicache/_0613_ ), .ZN(\myifu/myicache/_0882_ ) );
OAI211_X2 \myifu/myicache/_2327_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(fanout_net_24 ), .C2(\myifu/myicache/_0581_ ), .ZN(\myifu/myicache/_0883_ ) );
NOR2_X1 \myifu/myicache/_2328_ ( .A1(\myifu/myicache/_1063_ ), .A2(\myifu/myicache/_0517_ ), .ZN(\myifu/myicache/_0884_ ) );
OAI21_X1 \myifu/myicache/_2329_ ( .A(\myifu/myicache/_1034_ ), .B1(\myifu/myicache/_1038_ ), .B2(\myifu/myicache/_0549_ ), .ZN(\myifu/myicache/_0885_ ) );
OAI221_X1 \myifu/myicache/_2330_ ( .A(\myifu/myicache/_0881_ ), .B1(\myifu/myicache/_0882_ ), .B2(\myifu/myicache/_0883_ ), .C1(\myifu/myicache/_0884_ ), .C2(\myifu/myicache/_0885_ ), .ZN(\myifu/myicache/_0677_ ) );
MUX2_X1 \myifu/myicache/_2331_ ( .A(\myifu/myicache/_0391_ ), .B(\myifu/myicache/_0423_ ), .S(\myifu/myicache/_1063_ ), .Z(\myifu/myicache/_0886_ ) );
MUX2_X1 \myifu/myicache/_2332_ ( .A(\myifu/myicache/_0519_ ), .B(\myifu/myicache/_0551_ ), .S(\myifu/myicache/_1063_ ), .Z(\myifu/myicache/_0887_ ) );
AOI22_X1 \myifu/myicache/_2333_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0886_ ), .B1(\myifu/myicache/_0887_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0888_ ) );
NOR2_X1 \myifu/myicache/_2334_ ( .A1(\myifu/myicache/_1037_ ), .A2(\myifu/myicache/_0615_ ), .ZN(\myifu/myicache/_0889_ ) );
OAI211_X2 \myifu/myicache/_2335_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(\myifu/myicache/_1063_ ), .C2(\myifu/myicache/_0583_ ), .ZN(\myifu/myicache/_0890_ ) );
NOR2_X1 \myifu/myicache/_2336_ ( .A1(\myifu/myicache/_1043_ ), .A2(\myifu/myicache/_0487_ ), .ZN(\myifu/myicache/_0891_ ) );
OAI211_X2 \myifu/myicache/_2337_ ( .A(\myifu/myicache/_1040_ ), .B(\myifu/myicache/_0688_ ), .C1(\myifu/myicache/_1063_ ), .C2(\myifu/myicache/_0455_ ), .ZN(\myifu/myicache/_0892_ ) );
OAI221_X1 \myifu/myicache/_2338_ ( .A(\myifu/myicache/_0888_ ), .B1(\myifu/myicache/_0889_ ), .B2(\myifu/myicache/_0890_ ), .C1(\myifu/myicache/_0891_ ), .C2(\myifu/myicache/_0892_ ), .ZN(\myifu/myicache/_0679_ ) );
MUX2_X1 \myifu/myicache/_2339_ ( .A(\myifu/myicache/_0392_ ), .B(\myifu/myicache/_0424_ ), .S(\myifu/myicache/_1063_ ), .Z(\myifu/myicache/_0893_ ) );
MUX2_X1 \myifu/myicache/_2340_ ( .A(\myifu/myicache/_0520_ ), .B(\myifu/myicache/_0552_ ), .S(\myifu/myicache/_1063_ ), .Z(\myifu/myicache/_0894_ ) );
AOI22_X1 \myifu/myicache/_2341_ ( .A1(\myifu/myicache/_0815_ ), .A2(\myifu/myicache/_0893_ ), .B1(\myifu/myicache/_0894_ ), .B2(\myifu/myicache/_0794_ ), .ZN(\myifu/myicache/_0895_ ) );
NOR2_X1 \myifu/myicache/_2342_ ( .A1(\myifu/myicache/_1037_ ), .A2(\myifu/myicache/_0616_ ), .ZN(\myifu/myicache/_0896_ ) );
OAI211_X2 \myifu/myicache/_2343_ ( .A(\myifu/myicache/_0688_ ), .B(\myifu/myicache/_0689_ ), .C1(\myifu/myicache/_1063_ ), .C2(\myifu/myicache/_0584_ ), .ZN(\myifu/myicache/_0897_ ) );
NOR2_X1 \myifu/myicache/_2344_ ( .A1(\myifu/myicache/_1043_ ), .A2(\myifu/myicache/_0488_ ), .ZN(\myifu/myicache/_0898_ ) );
OAI211_X2 \myifu/myicache/_2345_ ( .A(\myifu/myicache/_1040_ ), .B(\myifu/myicache/_0688_ ), .C1(\myifu/myicache/_1063_ ), .C2(\myifu/myicache/_0456_ ), .ZN(\myifu/myicache/_0899_ ) );
OAI221_X1 \myifu/myicache/_2346_ ( .A(\myifu/myicache/_0895_ ), .B1(\myifu/myicache/_0896_ ), .B2(\myifu/myicache/_0897_ ), .C1(\myifu/myicache/_0898_ ), .C2(\myifu/myicache/_0899_ ), .ZN(\myifu/myicache/_0680_ ) );
INV_X32 \myifu/myicache/_2347_ ( .A(\myifu/myicache/_1064_ ), .ZN(\myifu/myicache/_0900_ ) );
AND2_X4 \myifu/myicache/_2348_ ( .A1(\myifu/myicache/_0900_ ), .A2(\myifu/myicache/_1233_ ), .ZN(\myifu/myicache/_0901_ ) );
AND2_X4 \myifu/myicache/_2349_ ( .A1(\myifu/myicache/_0901_ ), .A2(\myifu/myicache/_0960_ ), .ZN(\myifu/myicache/_0902_ ) );
NAND2_X4 \myifu/myicache/_2350_ ( .A1(\myifu/myicache/_0902_ ), .A2(\myifu/myicache/_1063_ ), .ZN(\myifu/myicache/_0903_ ) );
BUF_X4 \myifu/myicache/_2351_ ( .A(\myifu/myicache/_0903_ ), .Z(\myifu/myicache/_0904_ ) );
MUX2_X1 \myifu/myicache/_2352_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0528_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0000_ ) );
MUX2_X1 \myifu/myicache/_2353_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0539_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0001_ ) );
MUX2_X1 \myifu/myicache/_2354_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0550_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0002_ ) );
MUX2_X1 \myifu/myicache/_2355_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0553_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0003_ ) );
MUX2_X1 \myifu/myicache/_2356_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0554_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0004_ ) );
MUX2_X1 \myifu/myicache/_2357_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0555_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0005_ ) );
MUX2_X1 \myifu/myicache/_2358_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0556_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0006_ ) );
MUX2_X1 \myifu/myicache/_2359_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0557_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0007_ ) );
MUX2_X1 \myifu/myicache/_2360_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0558_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0008_ ) );
MUX2_X1 \myifu/myicache/_2361_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0559_ ), .S(\myifu/myicache/_0904_ ), .Z(\myifu/myicache/_0009_ ) );
BUF_X4 \myifu/myicache/_2362_ ( .A(\myifu/myicache/_0903_ ), .Z(\myifu/myicache/_0905_ ) );
MUX2_X1 \myifu/myicache/_2363_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0529_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0010_ ) );
MUX2_X1 \myifu/myicache/_2364_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0530_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0011_ ) );
MUX2_X1 \myifu/myicache/_2365_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0531_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0012_ ) );
MUX2_X1 \myifu/myicache/_2366_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0532_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0013_ ) );
MUX2_X1 \myifu/myicache/_2367_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0533_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0014_ ) );
MUX2_X1 \myifu/myicache/_2368_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0534_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0015_ ) );
MUX2_X1 \myifu/myicache/_2369_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0535_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0016_ ) );
MUX2_X1 \myifu/myicache/_2370_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0536_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0017_ ) );
MUX2_X1 \myifu/myicache/_2371_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0537_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0018_ ) );
MUX2_X1 \myifu/myicache/_2372_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0538_ ), .S(\myifu/myicache/_0905_ ), .Z(\myifu/myicache/_0019_ ) );
BUF_X4 \myifu/myicache/_2373_ ( .A(\myifu/myicache/_0903_ ), .Z(\myifu/myicache/_0906_ ) );
MUX2_X1 \myifu/myicache/_2374_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0540_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0020_ ) );
MUX2_X1 \myifu/myicache/_2375_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0541_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0021_ ) );
MUX2_X1 \myifu/myicache/_2376_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0542_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0022_ ) );
MUX2_X1 \myifu/myicache/_2377_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0543_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0023_ ) );
MUX2_X1 \myifu/myicache/_2378_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0544_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0024_ ) );
MUX2_X1 \myifu/myicache/_2379_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0545_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0025_ ) );
MUX2_X1 \myifu/myicache/_2380_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0546_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0026_ ) );
MUX2_X1 \myifu/myicache/_2381_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0547_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0027_ ) );
MUX2_X1 \myifu/myicache/_2382_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0548_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0028_ ) );
MUX2_X1 \myifu/myicache/_2383_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0549_ ), .S(\myifu/myicache/_0906_ ), .Z(\myifu/myicache/_0029_ ) );
MUX2_X1 \myifu/myicache/_2384_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0551_ ), .S(\myifu/myicache/_0903_ ), .Z(\myifu/myicache/_0030_ ) );
MUX2_X1 \myifu/myicache/_2385_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0552_ ), .S(\myifu/myicache/_0903_ ), .Z(\myifu/myicache/_0031_ ) );
NAND2_X4 \myifu/myicache/_2386_ ( .A1(\myifu/myicache/_0902_ ), .A2(\myifu/myicache/_1036_ ), .ZN(\myifu/myicache/_0907_ ) );
BUF_X4 \myifu/myicache/_2387_ ( .A(\myifu/myicache/_0907_ ), .Z(\myifu/myicache/_0908_ ) );
MUX2_X1 \myifu/myicache/_2388_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0496_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0032_ ) );
MUX2_X1 \myifu/myicache/_2389_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0507_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0033_ ) );
MUX2_X1 \myifu/myicache/_2390_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0518_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0034_ ) );
MUX2_X1 \myifu/myicache/_2391_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0521_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0035_ ) );
MUX2_X1 \myifu/myicache/_2392_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0522_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0036_ ) );
MUX2_X1 \myifu/myicache/_2393_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0523_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0037_ ) );
MUX2_X1 \myifu/myicache/_2394_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0524_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0038_ ) );
MUX2_X1 \myifu/myicache/_2395_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0525_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0039_ ) );
MUX2_X1 \myifu/myicache/_2396_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0526_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0040_ ) );
MUX2_X1 \myifu/myicache/_2397_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0527_ ), .S(\myifu/myicache/_0908_ ), .Z(\myifu/myicache/_0041_ ) );
BUF_X4 \myifu/myicache/_2398_ ( .A(\myifu/myicache/_0907_ ), .Z(\myifu/myicache/_0909_ ) );
MUX2_X1 \myifu/myicache/_2399_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0497_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0042_ ) );
MUX2_X1 \myifu/myicache/_2400_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0498_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0043_ ) );
MUX2_X1 \myifu/myicache/_2401_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0499_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0044_ ) );
MUX2_X1 \myifu/myicache/_2402_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0500_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0045_ ) );
MUX2_X1 \myifu/myicache/_2403_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0501_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0046_ ) );
MUX2_X1 \myifu/myicache/_2404_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0502_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0047_ ) );
MUX2_X1 \myifu/myicache/_2405_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0503_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0048_ ) );
MUX2_X1 \myifu/myicache/_2406_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0504_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0049_ ) );
MUX2_X1 \myifu/myicache/_2407_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0505_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0050_ ) );
MUX2_X1 \myifu/myicache/_2408_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0506_ ), .S(\myifu/myicache/_0909_ ), .Z(\myifu/myicache/_0051_ ) );
BUF_X4 \myifu/myicache/_2409_ ( .A(\myifu/myicache/_0907_ ), .Z(\myifu/myicache/_0910_ ) );
MUX2_X1 \myifu/myicache/_2410_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0508_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0052_ ) );
MUX2_X1 \myifu/myicache/_2411_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0509_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0053_ ) );
MUX2_X1 \myifu/myicache/_2412_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0510_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0054_ ) );
MUX2_X1 \myifu/myicache/_2413_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0511_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0055_ ) );
MUX2_X1 \myifu/myicache/_2414_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0512_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0056_ ) );
MUX2_X1 \myifu/myicache/_2415_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0513_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0057_ ) );
MUX2_X1 \myifu/myicache/_2416_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0514_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0058_ ) );
MUX2_X1 \myifu/myicache/_2417_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0515_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0059_ ) );
MUX2_X1 \myifu/myicache/_2418_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0516_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0060_ ) );
MUX2_X1 \myifu/myicache/_2419_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0517_ ), .S(\myifu/myicache/_0910_ ), .Z(\myifu/myicache/_0061_ ) );
MUX2_X1 \myifu/myicache/_2420_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0519_ ), .S(\myifu/myicache/_0907_ ), .Z(\myifu/myicache/_0062_ ) );
MUX2_X1 \myifu/myicache/_2421_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0520_ ), .S(\myifu/myicache/_0907_ ), .Z(\myifu/myicache/_0063_ ) );
AND2_X4 \myifu/myicache/_2422_ ( .A1(\myifu/myicache/_0901_ ), .A2(\myifu/myicache/_0971_ ), .ZN(\myifu/myicache/_0911_ ) );
BUF_X16 \myifu/myicache/_2423_ ( .A(\myifu/myicache/_0911_ ), .Z(\myifu/myicache/_0912_ ) );
NAND2_X4 \myifu/myicache/_2424_ ( .A1(\myifu/myicache/_0912_ ), .A2(\myifu/myicache/_1036_ ), .ZN(\myifu/myicache/_0913_ ) );
BUF_X8 \myifu/myicache/_2425_ ( .A(\myifu/myicache/_0913_ ), .Z(\myifu/myicache/_0914_ ) );
MUX2_X1 \myifu/myicache/_2426_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0560_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0064_ ) );
MUX2_X1 \myifu/myicache/_2427_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0571_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0065_ ) );
MUX2_X1 \myifu/myicache/_2428_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0582_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0066_ ) );
MUX2_X1 \myifu/myicache/_2429_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0585_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0067_ ) );
MUX2_X1 \myifu/myicache/_2430_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0586_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0068_ ) );
MUX2_X1 \myifu/myicache/_2431_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0587_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0069_ ) );
MUX2_X1 \myifu/myicache/_2432_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0588_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0070_ ) );
MUX2_X1 \myifu/myicache/_2433_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0589_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0071_ ) );
MUX2_X1 \myifu/myicache/_2434_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0590_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0072_ ) );
MUX2_X1 \myifu/myicache/_2435_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0591_ ), .S(\myifu/myicache/_0914_ ), .Z(\myifu/myicache/_0073_ ) );
BUF_X8 \myifu/myicache/_2436_ ( .A(\myifu/myicache/_0913_ ), .Z(\myifu/myicache/_0915_ ) );
MUX2_X1 \myifu/myicache/_2437_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0561_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0074_ ) );
MUX2_X1 \myifu/myicache/_2438_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0562_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0075_ ) );
MUX2_X1 \myifu/myicache/_2439_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0563_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0076_ ) );
MUX2_X1 \myifu/myicache/_2440_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0564_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0077_ ) );
MUX2_X1 \myifu/myicache/_2441_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0565_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0078_ ) );
MUX2_X1 \myifu/myicache/_2442_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0566_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0079_ ) );
MUX2_X1 \myifu/myicache/_2443_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0567_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0080_ ) );
MUX2_X1 \myifu/myicache/_2444_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0568_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0081_ ) );
MUX2_X1 \myifu/myicache/_2445_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0569_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0082_ ) );
MUX2_X1 \myifu/myicache/_2446_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0570_ ), .S(\myifu/myicache/_0915_ ), .Z(\myifu/myicache/_0083_ ) );
BUF_X8 \myifu/myicache/_2447_ ( .A(\myifu/myicache/_0913_ ), .Z(\myifu/myicache/_0916_ ) );
MUX2_X1 \myifu/myicache/_2448_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0572_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0084_ ) );
MUX2_X1 \myifu/myicache/_2449_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0573_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0085_ ) );
MUX2_X1 \myifu/myicache/_2450_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0574_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0086_ ) );
MUX2_X1 \myifu/myicache/_2451_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0575_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0087_ ) );
MUX2_X1 \myifu/myicache/_2452_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0576_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0088_ ) );
MUX2_X1 \myifu/myicache/_2453_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0577_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0089_ ) );
MUX2_X1 \myifu/myicache/_2454_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0578_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0090_ ) );
MUX2_X1 \myifu/myicache/_2455_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0579_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0091_ ) );
MUX2_X1 \myifu/myicache/_2456_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0580_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0092_ ) );
MUX2_X1 \myifu/myicache/_2457_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0581_ ), .S(\myifu/myicache/_0916_ ), .Z(\myifu/myicache/_0093_ ) );
MUX2_X1 \myifu/myicache/_2458_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0583_ ), .S(\myifu/myicache/_0913_ ), .Z(\myifu/myicache/_0094_ ) );
MUX2_X1 \myifu/myicache/_2459_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0584_ ), .S(\myifu/myicache/_0913_ ), .Z(\myifu/myicache/_0095_ ) );
AND2_X1 \myifu/myicache/_2460_ ( .A1(\myifu/myicache/_0900_ ), .A2(\myifu/myicache/_1229_ ), .ZN(\myifu/myicache/_0917_ ) );
BUF_X4 \myifu/myicache/_2461_ ( .A(\myifu/myicache/_0902_ ), .Z(\myifu/myicache/_0918_ ) );
BUF_X8 \myifu/myicache/_2462_ ( .A(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0919_ ) );
MUX2_X1 \myifu/myicache/_2463_ ( .A(\myifu/myicache/_0917_ ), .B(\myifu/myicache/_1231_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0096_ ) );
AND2_X1 \myifu/myicache/_2464_ ( .A1(\myifu/myicache/_0900_ ), .A2(\myifu/myicache/_1227_ ), .ZN(\myifu/myicache/_0920_ ) );
AND2_X4 \myifu/myicache/_2465_ ( .A1(\myifu/myicache/_0901_ ), .A2(\myifu/myicache/_0963_ ), .ZN(\myifu/myicache/_0921_ ) );
BUF_X4 \myifu/myicache/_2466_ ( .A(\myifu/myicache/_0921_ ), .Z(\myifu/myicache/_0922_ ) );
BUF_X4 \myifu/myicache/_2467_ ( .A(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0923_ ) );
MUX2_X1 \myifu/myicache/_2468_ ( .A(\myifu/myicache/_0920_ ), .B(\myifu/myicache/_1231_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0097_ ) );
AND2_X4 \myifu/myicache/_2469_ ( .A1(\myifu/myicache/_0958_ ), .A2(\myifu/myicache/_0901_ ), .ZN(\myifu/myicache/_0924_ ) );
NAND2_X4 \myifu/myicache/_2470_ ( .A1(\myifu/myicache/_0924_ ), .A2(\myifu/myicache/_1036_ ), .ZN(\myifu/myicache/_0925_ ) );
BUF_X4 \myifu/myicache/_2471_ ( .A(\myifu/myicache/_0925_ ), .Z(\myifu/myicache/_0926_ ) );
MUX2_X1 \myifu/myicache/_2472_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0432_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0098_ ) );
MUX2_X1 \myifu/myicache/_2473_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0443_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0099_ ) );
MUX2_X1 \myifu/myicache/_2474_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0454_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0100_ ) );
MUX2_X1 \myifu/myicache/_2475_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0457_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0101_ ) );
MUX2_X1 \myifu/myicache/_2476_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0458_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0102_ ) );
MUX2_X1 \myifu/myicache/_2477_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0459_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0103_ ) );
MUX2_X1 \myifu/myicache/_2478_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0460_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0104_ ) );
MUX2_X1 \myifu/myicache/_2479_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0461_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0105_ ) );
MUX2_X1 \myifu/myicache/_2480_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0462_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0106_ ) );
MUX2_X1 \myifu/myicache/_2481_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0463_ ), .S(\myifu/myicache/_0926_ ), .Z(\myifu/myicache/_0107_ ) );
BUF_X4 \myifu/myicache/_2482_ ( .A(\myifu/myicache/_0925_ ), .Z(\myifu/myicache/_0927_ ) );
MUX2_X1 \myifu/myicache/_2483_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0433_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0108_ ) );
MUX2_X1 \myifu/myicache/_2484_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0434_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0109_ ) );
MUX2_X1 \myifu/myicache/_2485_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0435_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0110_ ) );
MUX2_X1 \myifu/myicache/_2486_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0436_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0111_ ) );
MUX2_X1 \myifu/myicache/_2487_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0437_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0112_ ) );
MUX2_X1 \myifu/myicache/_2488_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0438_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0113_ ) );
MUX2_X1 \myifu/myicache/_2489_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0439_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0114_ ) );
MUX2_X1 \myifu/myicache/_2490_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0440_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0115_ ) );
MUX2_X1 \myifu/myicache/_2491_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0441_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0116_ ) );
MUX2_X1 \myifu/myicache/_2492_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0442_ ), .S(\myifu/myicache/_0927_ ), .Z(\myifu/myicache/_0117_ ) );
BUF_X4 \myifu/myicache/_2493_ ( .A(\myifu/myicache/_0925_ ), .Z(\myifu/myicache/_0928_ ) );
MUX2_X1 \myifu/myicache/_2494_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0444_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0118_ ) );
MUX2_X1 \myifu/myicache/_2495_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0445_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0119_ ) );
MUX2_X1 \myifu/myicache/_2496_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0446_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0120_ ) );
MUX2_X1 \myifu/myicache/_2497_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0447_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0121_ ) );
MUX2_X1 \myifu/myicache/_2498_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0448_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0122_ ) );
MUX2_X1 \myifu/myicache/_2499_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0449_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0123_ ) );
MUX2_X1 \myifu/myicache/_2500_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0450_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0124_ ) );
MUX2_X1 \myifu/myicache/_2501_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0451_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0125_ ) );
MUX2_X1 \myifu/myicache/_2502_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0452_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0126_ ) );
MUX2_X1 \myifu/myicache/_2503_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0453_ ), .S(\myifu/myicache/_0928_ ), .Z(\myifu/myicache/_0127_ ) );
MUX2_X1 \myifu/myicache/_2504_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0455_ ), .S(\myifu/myicache/_0925_ ), .Z(\myifu/myicache/_0128_ ) );
MUX2_X1 \myifu/myicache/_2505_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0456_ ), .S(\myifu/myicache/_0925_ ), .Z(\myifu/myicache/_0129_ ) );
NAND2_X4 \myifu/myicache/_2506_ ( .A1(\myifu/myicache/_0921_ ), .A2(\myifu/myicache/_1063_ ), .ZN(\myifu/myicache/_0929_ ) );
BUF_X4 \myifu/myicache/_2507_ ( .A(\myifu/myicache/_0929_ ), .Z(\myifu/myicache/_0930_ ) );
MUX2_X1 \myifu/myicache/_2508_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0400_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0130_ ) );
MUX2_X1 \myifu/myicache/_2509_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0411_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0131_ ) );
MUX2_X1 \myifu/myicache/_2510_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0422_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0132_ ) );
MUX2_X1 \myifu/myicache/_2511_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0425_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0133_ ) );
MUX2_X1 \myifu/myicache/_2512_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0426_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0134_ ) );
MUX2_X1 \myifu/myicache/_2513_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0427_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0135_ ) );
MUX2_X1 \myifu/myicache/_2514_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0428_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0136_ ) );
MUX2_X1 \myifu/myicache/_2515_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0429_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0137_ ) );
MUX2_X1 \myifu/myicache/_2516_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0430_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0138_ ) );
MUX2_X1 \myifu/myicache/_2517_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0431_ ), .S(\myifu/myicache/_0930_ ), .Z(\myifu/myicache/_0139_ ) );
BUF_X4 \myifu/myicache/_2518_ ( .A(\myifu/myicache/_0929_ ), .Z(\myifu/myicache/_0931_ ) );
MUX2_X1 \myifu/myicache/_2519_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0401_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0140_ ) );
MUX2_X1 \myifu/myicache/_2520_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0402_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0141_ ) );
MUX2_X1 \myifu/myicache/_2521_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0403_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0142_ ) );
MUX2_X1 \myifu/myicache/_2522_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0404_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0143_ ) );
MUX2_X1 \myifu/myicache/_2523_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0405_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0144_ ) );
MUX2_X1 \myifu/myicache/_2524_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0406_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0145_ ) );
MUX2_X1 \myifu/myicache/_2525_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0407_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0146_ ) );
MUX2_X1 \myifu/myicache/_2526_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0408_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0147_ ) );
MUX2_X1 \myifu/myicache/_2527_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0409_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0148_ ) );
MUX2_X1 \myifu/myicache/_2528_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0410_ ), .S(\myifu/myicache/_0931_ ), .Z(\myifu/myicache/_0149_ ) );
BUF_X4 \myifu/myicache/_2529_ ( .A(\myifu/myicache/_0929_ ), .Z(\myifu/myicache/_0932_ ) );
MUX2_X1 \myifu/myicache/_2530_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0412_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0150_ ) );
MUX2_X1 \myifu/myicache/_2531_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0413_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0151_ ) );
MUX2_X1 \myifu/myicache/_2532_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0414_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0152_ ) );
MUX2_X1 \myifu/myicache/_2533_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0415_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0153_ ) );
MUX2_X1 \myifu/myicache/_2534_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0416_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0154_ ) );
MUX2_X1 \myifu/myicache/_2535_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0417_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0155_ ) );
MUX2_X1 \myifu/myicache/_2536_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0418_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0156_ ) );
MUX2_X1 \myifu/myicache/_2537_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0419_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0157_ ) );
MUX2_X1 \myifu/myicache/_2538_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0420_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0158_ ) );
MUX2_X1 \myifu/myicache/_2539_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0421_ ), .S(\myifu/myicache/_0932_ ), .Z(\myifu/myicache/_0159_ ) );
MUX2_X1 \myifu/myicache/_2540_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0423_ ), .S(\myifu/myicache/_0929_ ), .Z(\myifu/myicache/_0160_ ) );
MUX2_X1 \myifu/myicache/_2541_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0424_ ), .S(\myifu/myicache/_0929_ ), .Z(\myifu/myicache/_0161_ ) );
NAND2_X4 \myifu/myicache/_2542_ ( .A1(\myifu/myicache/_0921_ ), .A2(\myifu/myicache/_1036_ ), .ZN(\myifu/myicache/_0933_ ) );
BUF_X4 \myifu/myicache/_2543_ ( .A(\myifu/myicache/_0933_ ), .Z(\myifu/myicache/_0934_ ) );
MUX2_X1 \myifu/myicache/_2544_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0368_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0162_ ) );
MUX2_X1 \myifu/myicache/_2545_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0379_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0163_ ) );
MUX2_X1 \myifu/myicache/_2546_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0390_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0164_ ) );
MUX2_X1 \myifu/myicache/_2547_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0393_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0165_ ) );
MUX2_X1 \myifu/myicache/_2548_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0394_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0166_ ) );
MUX2_X1 \myifu/myicache/_2549_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0395_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0167_ ) );
MUX2_X1 \myifu/myicache/_2550_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0396_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0168_ ) );
MUX2_X1 \myifu/myicache/_2551_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0397_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0169_ ) );
MUX2_X1 \myifu/myicache/_2552_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0398_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0170_ ) );
MUX2_X1 \myifu/myicache/_2553_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0399_ ), .S(\myifu/myicache/_0934_ ), .Z(\myifu/myicache/_0171_ ) );
BUF_X4 \myifu/myicache/_2554_ ( .A(\myifu/myicache/_0933_ ), .Z(\myifu/myicache/_0935_ ) );
MUX2_X1 \myifu/myicache/_2555_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0369_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0172_ ) );
MUX2_X1 \myifu/myicache/_2556_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0370_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0173_ ) );
MUX2_X1 \myifu/myicache/_2557_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0371_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0174_ ) );
MUX2_X1 \myifu/myicache/_2558_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0372_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0175_ ) );
MUX2_X1 \myifu/myicache/_2559_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0373_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0176_ ) );
MUX2_X1 \myifu/myicache/_2560_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0374_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0177_ ) );
MUX2_X1 \myifu/myicache/_2561_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0375_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0178_ ) );
MUX2_X1 \myifu/myicache/_2562_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0376_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0179_ ) );
MUX2_X1 \myifu/myicache/_2563_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0377_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0180_ ) );
MUX2_X1 \myifu/myicache/_2564_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0378_ ), .S(\myifu/myicache/_0935_ ), .Z(\myifu/myicache/_0181_ ) );
BUF_X4 \myifu/myicache/_2565_ ( .A(\myifu/myicache/_0933_ ), .Z(\myifu/myicache/_0936_ ) );
MUX2_X1 \myifu/myicache/_2566_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0380_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0182_ ) );
MUX2_X1 \myifu/myicache/_2567_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0381_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0183_ ) );
MUX2_X1 \myifu/myicache/_2568_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0382_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0184_ ) );
MUX2_X1 \myifu/myicache/_2569_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0383_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0185_ ) );
MUX2_X1 \myifu/myicache/_2570_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0384_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0186_ ) );
MUX2_X1 \myifu/myicache/_2571_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0385_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0187_ ) );
MUX2_X1 \myifu/myicache/_2572_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0386_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0188_ ) );
MUX2_X1 \myifu/myicache/_2573_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0387_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0189_ ) );
MUX2_X1 \myifu/myicache/_2574_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0388_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0190_ ) );
MUX2_X1 \myifu/myicache/_2575_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0389_ ), .S(\myifu/myicache/_0936_ ), .Z(\myifu/myicache/_0191_ ) );
MUX2_X1 \myifu/myicache/_2576_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0391_ ), .S(\myifu/myicache/_0933_ ), .Z(\myifu/myicache/_0192_ ) );
MUX2_X1 \myifu/myicache/_2577_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0392_ ), .S(\myifu/myicache/_0933_ ), .Z(\myifu/myicache/_0193_ ) );
NAND4_X1 \myifu/myicache/_2578_ ( .A1(\myifu/myicache/_0972_ ), .A2(\myifu/myicache/_0900_ ), .A3(\myifu/myicache/_1233_ ), .A4(\myifu/myicache/_1231_ ), .ZN(\myifu/myicache/_0937_ ) );
NAND3_X1 \myifu/myicache/_2579_ ( .A1(\myifu/myicache/_0688_ ), .A2(\myifu/myicache/_0689_ ), .A3(\myifu/myicache/_1233_ ), .ZN(\myifu/myicache/_0938_ ) );
NAND3_X1 \myifu/myicache/_2580_ ( .A1(\myifu/myicache/_0938_ ), .A2(\myifu/myicache/_0900_ ), .A3(\myifu/myicache/_1230_ ), .ZN(\myifu/myicache/_0939_ ) );
NAND2_X1 \myifu/myicache/_2581_ ( .A1(\myifu/myicache/_0937_ ), .A2(\myifu/myicache/_0939_ ), .ZN(\myifu/myicache/_0194_ ) );
NAND2_X4 \myifu/myicache/_2582_ ( .A1(\myifu/myicache/_0924_ ), .A2(\myifu/myicache/_1063_ ), .ZN(\myifu/myicache/_0940_ ) );
BUF_X4 \myifu/myicache/_2583_ ( .A(\myifu/myicache/_0940_ ), .Z(\myifu/myicache/_0941_ ) );
MUX2_X1 \myifu/myicache/_2584_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0464_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0195_ ) );
MUX2_X1 \myifu/myicache/_2585_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0475_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0196_ ) );
MUX2_X1 \myifu/myicache/_2586_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0486_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0197_ ) );
MUX2_X1 \myifu/myicache/_2587_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0489_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0198_ ) );
MUX2_X1 \myifu/myicache/_2588_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0490_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0199_ ) );
MUX2_X1 \myifu/myicache/_2589_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0491_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0200_ ) );
MUX2_X1 \myifu/myicache/_2590_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0492_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0201_ ) );
MUX2_X1 \myifu/myicache/_2591_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0493_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0202_ ) );
MUX2_X1 \myifu/myicache/_2592_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0494_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0203_ ) );
MUX2_X1 \myifu/myicache/_2593_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0495_ ), .S(\myifu/myicache/_0941_ ), .Z(\myifu/myicache/_0204_ ) );
BUF_X4 \myifu/myicache/_2594_ ( .A(\myifu/myicache/_0940_ ), .Z(\myifu/myicache/_0942_ ) );
MUX2_X1 \myifu/myicache/_2595_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0465_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0205_ ) );
MUX2_X1 \myifu/myicache/_2596_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0466_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0206_ ) );
MUX2_X1 \myifu/myicache/_2597_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0467_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0207_ ) );
MUX2_X1 \myifu/myicache/_2598_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0468_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0208_ ) );
MUX2_X1 \myifu/myicache/_2599_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0469_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0209_ ) );
MUX2_X1 \myifu/myicache/_2600_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0470_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0210_ ) );
MUX2_X1 \myifu/myicache/_2601_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0471_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0211_ ) );
MUX2_X1 \myifu/myicache/_2602_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0472_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0212_ ) );
MUX2_X1 \myifu/myicache/_2603_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0473_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0213_ ) );
MUX2_X1 \myifu/myicache/_2604_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0474_ ), .S(\myifu/myicache/_0942_ ), .Z(\myifu/myicache/_0214_ ) );
BUF_X4 \myifu/myicache/_2605_ ( .A(\myifu/myicache/_0940_ ), .Z(\myifu/myicache/_0943_ ) );
MUX2_X1 \myifu/myicache/_2606_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0476_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0215_ ) );
MUX2_X1 \myifu/myicache/_2607_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0477_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0216_ ) );
MUX2_X1 \myifu/myicache/_2608_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0478_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0217_ ) );
MUX2_X1 \myifu/myicache/_2609_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0479_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0218_ ) );
MUX2_X1 \myifu/myicache/_2610_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0480_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0219_ ) );
MUX2_X1 \myifu/myicache/_2611_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0481_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0220_ ) );
MUX2_X1 \myifu/myicache/_2612_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0482_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0221_ ) );
MUX2_X1 \myifu/myicache/_2613_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0483_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0222_ ) );
MUX2_X1 \myifu/myicache/_2614_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0484_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0223_ ) );
MUX2_X1 \myifu/myicache/_2615_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0485_ ), .S(\myifu/myicache/_0943_ ), .Z(\myifu/myicache/_0224_ ) );
MUX2_X1 \myifu/myicache/_2616_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0487_ ), .S(\myifu/myicache/_0940_ ), .Z(\myifu/myicache/_0225_ ) );
MUX2_X1 \myifu/myicache/_2617_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0488_ ), .S(\myifu/myicache/_0940_ ), .Z(\myifu/myicache/_0226_ ) );
MUX2_X1 \myifu/myicache/_2618_ ( .A(\myifu/myicache/_1119_ ), .B(\myifu/myicache/_1173_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0227_ ) );
MUX2_X1 \myifu/myicache/_2619_ ( .A(\myifu/myicache/_1130_ ), .B(\myifu/myicache/_1184_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0228_ ) );
MUX2_X1 \myifu/myicache/_2620_ ( .A(\myifu/myicache/_1138_ ), .B(\myifu/myicache/_1192_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0229_ ) );
MUX2_X1 \myifu/myicache/_2621_ ( .A(\myifu/myicache/_1139_ ), .B(\myifu/myicache/_1193_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0230_ ) );
MUX2_X1 \myifu/myicache/_2622_ ( .A(\myifu/myicache/_1140_ ), .B(\myifu/myicache/_1194_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0231_ ) );
MUX2_X1 \myifu/myicache/_2623_ ( .A(\myifu/myicache/_1141_ ), .B(\myifu/myicache/_1195_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0232_ ) );
MUX2_X1 \myifu/myicache/_2624_ ( .A(\myifu/myicache/_1142_ ), .B(\myifu/myicache/_1196_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0233_ ) );
MUX2_X1 \myifu/myicache/_2625_ ( .A(\myifu/myicache/_1143_ ), .B(\myifu/myicache/_1197_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0234_ ) );
MUX2_X1 \myifu/myicache/_2626_ ( .A(\myifu/myicache/_1144_ ), .B(\myifu/myicache/_1198_ ), .S(\myifu/myicache/_0919_ ), .Z(\myifu/myicache/_0235_ ) );
BUF_X4 \myifu/myicache/_2627_ ( .A(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0944_ ) );
MUX2_X1 \myifu/myicache/_2628_ ( .A(\myifu/myicache/_1145_ ), .B(\myifu/myicache/_1199_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0236_ ) );
MUX2_X1 \myifu/myicache/_2629_ ( .A(\myifu/myicache/_1120_ ), .B(\myifu/myicache/_1174_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0237_ ) );
MUX2_X1 \myifu/myicache/_2630_ ( .A(\myifu/myicache/_1121_ ), .B(\myifu/myicache/_1175_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0238_ ) );
MUX2_X1 \myifu/myicache/_2631_ ( .A(\myifu/myicache/_1122_ ), .B(\myifu/myicache/_1176_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0239_ ) );
MUX2_X1 \myifu/myicache/_2632_ ( .A(\myifu/myicache/_1123_ ), .B(\myifu/myicache/_1177_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0240_ ) );
MUX2_X1 \myifu/myicache/_2633_ ( .A(\myifu/myicache/_1124_ ), .B(\myifu/myicache/_1178_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0241_ ) );
MUX2_X1 \myifu/myicache/_2634_ ( .A(\myifu/myicache/_1125_ ), .B(\myifu/myicache/_1179_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0242_ ) );
MUX2_X1 \myifu/myicache/_2635_ ( .A(\myifu/myicache/_1126_ ), .B(\myifu/myicache/_1180_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0243_ ) );
MUX2_X1 \myifu/myicache/_2636_ ( .A(\myifu/myicache/_1127_ ), .B(\myifu/myicache/_1181_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0244_ ) );
MUX2_X1 \myifu/myicache/_2637_ ( .A(\myifu/myicache/_1128_ ), .B(\myifu/myicache/_1182_ ), .S(\myifu/myicache/_0944_ ), .Z(\myifu/myicache/_0245_ ) );
MUX2_X1 \myifu/myicache/_2638_ ( .A(\myifu/myicache/_1129_ ), .B(\myifu/myicache/_1183_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0246_ ) );
MUX2_X1 \myifu/myicache/_2639_ ( .A(\myifu/myicache/_1131_ ), .B(\myifu/myicache/_1185_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0247_ ) );
MUX2_X1 \myifu/myicache/_2640_ ( .A(\myifu/myicache/_1132_ ), .B(\myifu/myicache/_1186_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0248_ ) );
MUX2_X1 \myifu/myicache/_2641_ ( .A(\myifu/myicache/_1133_ ), .B(\myifu/myicache/_1187_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0249_ ) );
MUX2_X1 \myifu/myicache/_2642_ ( .A(\myifu/myicache/_1134_ ), .B(\myifu/myicache/_1188_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0250_ ) );
MUX2_X1 \myifu/myicache/_2643_ ( .A(\myifu/myicache/_1135_ ), .B(\myifu/myicache/_1189_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0251_ ) );
MUX2_X1 \myifu/myicache/_2644_ ( .A(\myifu/myicache/_1136_ ), .B(\myifu/myicache/_1190_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0252_ ) );
MUX2_X1 \myifu/myicache/_2645_ ( .A(\myifu/myicache/_1137_ ), .B(\myifu/myicache/_1191_ ), .S(\myifu/myicache/_0918_ ), .Z(\myifu/myicache/_0253_ ) );
BUF_X4 \myifu/myicache/_2646_ ( .A(\myifu/myicache/_0924_ ), .Z(\myifu/myicache/_0945_ ) );
BUF_X4 \myifu/myicache/_2647_ ( .A(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0946_ ) );
MUX2_X1 \myifu/myicache/_2648_ ( .A(\myifu/myicache/_1092_ ), .B(\myifu/myicache/_1173_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0254_ ) );
MUX2_X1 \myifu/myicache/_2649_ ( .A(\myifu/myicache/_1103_ ), .B(\myifu/myicache/_1184_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0255_ ) );
MUX2_X1 \myifu/myicache/_2650_ ( .A(\myifu/myicache/_1111_ ), .B(\myifu/myicache/_1192_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0256_ ) );
MUX2_X1 \myifu/myicache/_2651_ ( .A(\myifu/myicache/_1112_ ), .B(\myifu/myicache/_1193_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0257_ ) );
MUX2_X1 \myifu/myicache/_2652_ ( .A(\myifu/myicache/_1113_ ), .B(\myifu/myicache/_1194_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0258_ ) );
MUX2_X1 \myifu/myicache/_2653_ ( .A(\myifu/myicache/_1114_ ), .B(\myifu/myicache/_1195_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0259_ ) );
MUX2_X1 \myifu/myicache/_2654_ ( .A(\myifu/myicache/_1115_ ), .B(\myifu/myicache/_1196_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0260_ ) );
MUX2_X1 \myifu/myicache/_2655_ ( .A(\myifu/myicache/_1116_ ), .B(\myifu/myicache/_1197_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0261_ ) );
MUX2_X1 \myifu/myicache/_2656_ ( .A(\myifu/myicache/_1117_ ), .B(\myifu/myicache/_1198_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0262_ ) );
MUX2_X1 \myifu/myicache/_2657_ ( .A(\myifu/myicache/_1118_ ), .B(\myifu/myicache/_1199_ ), .S(\myifu/myicache/_0946_ ), .Z(\myifu/myicache/_0263_ ) );
BUF_X4 \myifu/myicache/_2658_ ( .A(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0947_ ) );
MUX2_X1 \myifu/myicache/_2659_ ( .A(\myifu/myicache/_1093_ ), .B(\myifu/myicache/_1174_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0264_ ) );
MUX2_X1 \myifu/myicache/_2660_ ( .A(\myifu/myicache/_1094_ ), .B(\myifu/myicache/_1175_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0265_ ) );
MUX2_X1 \myifu/myicache/_2661_ ( .A(\myifu/myicache/_1095_ ), .B(\myifu/myicache/_1176_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0266_ ) );
MUX2_X1 \myifu/myicache/_2662_ ( .A(\myifu/myicache/_1096_ ), .B(\myifu/myicache/_1177_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0267_ ) );
MUX2_X1 \myifu/myicache/_2663_ ( .A(\myifu/myicache/_1097_ ), .B(\myifu/myicache/_1178_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0268_ ) );
MUX2_X1 \myifu/myicache/_2664_ ( .A(\myifu/myicache/_1098_ ), .B(\myifu/myicache/_1179_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0269_ ) );
MUX2_X1 \myifu/myicache/_2665_ ( .A(\myifu/myicache/_1099_ ), .B(\myifu/myicache/_1180_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0270_ ) );
MUX2_X1 \myifu/myicache/_2666_ ( .A(\myifu/myicache/_1100_ ), .B(\myifu/myicache/_1181_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0271_ ) );
MUX2_X1 \myifu/myicache/_2667_ ( .A(\myifu/myicache/_1101_ ), .B(\myifu/myicache/_1182_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0272_ ) );
MUX2_X1 \myifu/myicache/_2668_ ( .A(\myifu/myicache/_1102_ ), .B(\myifu/myicache/_1183_ ), .S(\myifu/myicache/_0947_ ), .Z(\myifu/myicache/_0273_ ) );
MUX2_X1 \myifu/myicache/_2669_ ( .A(\myifu/myicache/_1104_ ), .B(\myifu/myicache/_1185_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0274_ ) );
MUX2_X1 \myifu/myicache/_2670_ ( .A(\myifu/myicache/_1105_ ), .B(\myifu/myicache/_1186_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0275_ ) );
MUX2_X1 \myifu/myicache/_2671_ ( .A(\myifu/myicache/_1106_ ), .B(\myifu/myicache/_1187_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0276_ ) );
MUX2_X1 \myifu/myicache/_2672_ ( .A(\myifu/myicache/_1107_ ), .B(\myifu/myicache/_1188_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0277_ ) );
MUX2_X1 \myifu/myicache/_2673_ ( .A(\myifu/myicache/_1108_ ), .B(\myifu/myicache/_1189_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0278_ ) );
MUX2_X1 \myifu/myicache/_2674_ ( .A(\myifu/myicache/_1109_ ), .B(\myifu/myicache/_1190_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0279_ ) );
MUX2_X1 \myifu/myicache/_2675_ ( .A(\myifu/myicache/_1110_ ), .B(\myifu/myicache/_1191_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0280_ ) );
MUX2_X1 \myifu/myicache/_2676_ ( .A(\myifu/myicache/_1065_ ), .B(\myifu/myicache/_1173_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0281_ ) );
MUX2_X1 \myifu/myicache/_2677_ ( .A(\myifu/myicache/_1076_ ), .B(\myifu/myicache/_1184_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0282_ ) );
MUX2_X1 \myifu/myicache/_2678_ ( .A(\myifu/myicache/_1084_ ), .B(\myifu/myicache/_1192_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0283_ ) );
MUX2_X1 \myifu/myicache/_2679_ ( .A(\myifu/myicache/_1085_ ), .B(\myifu/myicache/_1193_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0284_ ) );
MUX2_X1 \myifu/myicache/_2680_ ( .A(\myifu/myicache/_1086_ ), .B(\myifu/myicache/_1194_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0285_ ) );
MUX2_X1 \myifu/myicache/_2681_ ( .A(\myifu/myicache/_1087_ ), .B(\myifu/myicache/_1195_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0286_ ) );
MUX2_X1 \myifu/myicache/_2682_ ( .A(\myifu/myicache/_1088_ ), .B(\myifu/myicache/_1196_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0287_ ) );
MUX2_X1 \myifu/myicache/_2683_ ( .A(\myifu/myicache/_1089_ ), .B(\myifu/myicache/_1197_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0288_ ) );
MUX2_X1 \myifu/myicache/_2684_ ( .A(\myifu/myicache/_1090_ ), .B(\myifu/myicache/_1198_ ), .S(\myifu/myicache/_0923_ ), .Z(\myifu/myicache/_0289_ ) );
BUF_X8 \myifu/myicache/_2685_ ( .A(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0948_ ) );
MUX2_X1 \myifu/myicache/_2686_ ( .A(\myifu/myicache/_1091_ ), .B(\myifu/myicache/_1199_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0290_ ) );
MUX2_X1 \myifu/myicache/_2687_ ( .A(\myifu/myicache/_1066_ ), .B(\myifu/myicache/_1174_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0291_ ) );
MUX2_X1 \myifu/myicache/_2688_ ( .A(\myifu/myicache/_1067_ ), .B(\myifu/myicache/_1175_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0292_ ) );
MUX2_X1 \myifu/myicache/_2689_ ( .A(\myifu/myicache/_1068_ ), .B(\myifu/myicache/_1176_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0293_ ) );
MUX2_X1 \myifu/myicache/_2690_ ( .A(\myifu/myicache/_1069_ ), .B(\myifu/myicache/_1177_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0294_ ) );
MUX2_X1 \myifu/myicache/_2691_ ( .A(\myifu/myicache/_1070_ ), .B(\myifu/myicache/_1178_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0295_ ) );
MUX2_X1 \myifu/myicache/_2692_ ( .A(\myifu/myicache/_1071_ ), .B(\myifu/myicache/_1179_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0296_ ) );
MUX2_X1 \myifu/myicache/_2693_ ( .A(\myifu/myicache/_1072_ ), .B(\myifu/myicache/_1180_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0297_ ) );
MUX2_X1 \myifu/myicache/_2694_ ( .A(\myifu/myicache/_1073_ ), .B(\myifu/myicache/_1181_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0298_ ) );
MUX2_X1 \myifu/myicache/_2695_ ( .A(\myifu/myicache/_1074_ ), .B(\myifu/myicache/_1182_ ), .S(\myifu/myicache/_0948_ ), .Z(\myifu/myicache/_0299_ ) );
MUX2_X1 \myifu/myicache/_2696_ ( .A(\myifu/myicache/_1075_ ), .B(\myifu/myicache/_1183_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0300_ ) );
MUX2_X1 \myifu/myicache/_2697_ ( .A(\myifu/myicache/_1077_ ), .B(\myifu/myicache/_1185_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0301_ ) );
MUX2_X1 \myifu/myicache/_2698_ ( .A(\myifu/myicache/_1078_ ), .B(\myifu/myicache/_1186_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0302_ ) );
MUX2_X1 \myifu/myicache/_2699_ ( .A(\myifu/myicache/_1079_ ), .B(\myifu/myicache/_1187_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0303_ ) );
MUX2_X1 \myifu/myicache/_2700_ ( .A(\myifu/myicache/_1080_ ), .B(\myifu/myicache/_1188_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0304_ ) );
MUX2_X1 \myifu/myicache/_2701_ ( .A(\myifu/myicache/_1081_ ), .B(\myifu/myicache/_1189_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0305_ ) );
MUX2_X1 \myifu/myicache/_2702_ ( .A(\myifu/myicache/_1082_ ), .B(\myifu/myicache/_1190_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0306_ ) );
MUX2_X1 \myifu/myicache/_2703_ ( .A(\myifu/myicache/_1083_ ), .B(\myifu/myicache/_1191_ ), .S(\myifu/myicache/_0922_ ), .Z(\myifu/myicache/_0307_ ) );
NAND2_X4 \myifu/myicache/_2704_ ( .A1(\myifu/myicache/_0911_ ), .A2(\myifu/myicache/_1063_ ), .ZN(\myifu/myicache/_0949_ ) );
BUF_X4 \myifu/myicache/_2705_ ( .A(\myifu/myicache/_0949_ ), .Z(\myifu/myicache/_0950_ ) );
MUX2_X1 \myifu/myicache/_2706_ ( .A(\myifu/myicache/_0624_ ), .B(\myifu/myicache/_0592_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0308_ ) );
MUX2_X1 \myifu/myicache/_2707_ ( .A(\myifu/myicache/_0635_ ), .B(\myifu/myicache/_0603_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0309_ ) );
MUX2_X1 \myifu/myicache/_2708_ ( .A(\myifu/myicache/_0646_ ), .B(\myifu/myicache/_0614_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0310_ ) );
MUX2_X1 \myifu/myicache/_2709_ ( .A(\myifu/myicache/_0649_ ), .B(\myifu/myicache/_0617_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0311_ ) );
MUX2_X1 \myifu/myicache/_2710_ ( .A(\myifu/myicache/_0650_ ), .B(\myifu/myicache/_0618_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0312_ ) );
MUX2_X1 \myifu/myicache/_2711_ ( .A(\myifu/myicache/_0651_ ), .B(\myifu/myicache/_0619_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0313_ ) );
MUX2_X1 \myifu/myicache/_2712_ ( .A(\myifu/myicache/_0652_ ), .B(\myifu/myicache/_0620_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0314_ ) );
MUX2_X1 \myifu/myicache/_2713_ ( .A(\myifu/myicache/_0653_ ), .B(\myifu/myicache/_0621_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0315_ ) );
MUX2_X1 \myifu/myicache/_2714_ ( .A(\myifu/myicache/_0654_ ), .B(\myifu/myicache/_0622_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0316_ ) );
MUX2_X1 \myifu/myicache/_2715_ ( .A(\myifu/myicache/_0655_ ), .B(\myifu/myicache/_0623_ ), .S(\myifu/myicache/_0950_ ), .Z(\myifu/myicache/_0317_ ) );
BUF_X4 \myifu/myicache/_2716_ ( .A(\myifu/myicache/_0949_ ), .Z(\myifu/myicache/_0951_ ) );
MUX2_X1 \myifu/myicache/_2717_ ( .A(\myifu/myicache/_0625_ ), .B(\myifu/myicache/_0593_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0318_ ) );
MUX2_X1 \myifu/myicache/_2718_ ( .A(\myifu/myicache/_0626_ ), .B(\myifu/myicache/_0594_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0319_ ) );
MUX2_X1 \myifu/myicache/_2719_ ( .A(\myifu/myicache/_0627_ ), .B(\myifu/myicache/_0595_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0320_ ) );
MUX2_X1 \myifu/myicache/_2720_ ( .A(\myifu/myicache/_0628_ ), .B(\myifu/myicache/_0596_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0321_ ) );
MUX2_X1 \myifu/myicache/_2721_ ( .A(\myifu/myicache/_0629_ ), .B(\myifu/myicache/_0597_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0322_ ) );
MUX2_X1 \myifu/myicache/_2722_ ( .A(\myifu/myicache/_0630_ ), .B(\myifu/myicache/_0598_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0323_ ) );
MUX2_X1 \myifu/myicache/_2723_ ( .A(\myifu/myicache/_0631_ ), .B(\myifu/myicache/_0599_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0324_ ) );
MUX2_X1 \myifu/myicache/_2724_ ( .A(\myifu/myicache/_0632_ ), .B(\myifu/myicache/_0600_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0325_ ) );
MUX2_X1 \myifu/myicache/_2725_ ( .A(\myifu/myicache/_0633_ ), .B(\myifu/myicache/_0601_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0326_ ) );
MUX2_X1 \myifu/myicache/_2726_ ( .A(\myifu/myicache/_0634_ ), .B(\myifu/myicache/_0602_ ), .S(\myifu/myicache/_0951_ ), .Z(\myifu/myicache/_0327_ ) );
BUF_X4 \myifu/myicache/_2727_ ( .A(\myifu/myicache/_0949_ ), .Z(\myifu/myicache/_0952_ ) );
MUX2_X1 \myifu/myicache/_2728_ ( .A(\myifu/myicache/_0636_ ), .B(\myifu/myicache/_0604_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0328_ ) );
MUX2_X1 \myifu/myicache/_2729_ ( .A(\myifu/myicache/_0637_ ), .B(\myifu/myicache/_0605_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0329_ ) );
MUX2_X1 \myifu/myicache/_2730_ ( .A(\myifu/myicache/_0638_ ), .B(\myifu/myicache/_0606_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0330_ ) );
MUX2_X1 \myifu/myicache/_2731_ ( .A(\myifu/myicache/_0639_ ), .B(\myifu/myicache/_0607_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0331_ ) );
MUX2_X1 \myifu/myicache/_2732_ ( .A(\myifu/myicache/_0640_ ), .B(\myifu/myicache/_0608_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0332_ ) );
MUX2_X1 \myifu/myicache/_2733_ ( .A(\myifu/myicache/_0641_ ), .B(\myifu/myicache/_0609_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0333_ ) );
MUX2_X1 \myifu/myicache/_2734_ ( .A(\myifu/myicache/_0642_ ), .B(\myifu/myicache/_0610_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0334_ ) );
MUX2_X1 \myifu/myicache/_2735_ ( .A(\myifu/myicache/_0643_ ), .B(\myifu/myicache/_0611_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0335_ ) );
MUX2_X1 \myifu/myicache/_2736_ ( .A(\myifu/myicache/_0644_ ), .B(\myifu/myicache/_0612_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0336_ ) );
MUX2_X1 \myifu/myicache/_2737_ ( .A(\myifu/myicache/_0645_ ), .B(\myifu/myicache/_0613_ ), .S(\myifu/myicache/_0952_ ), .Z(\myifu/myicache/_0337_ ) );
MUX2_X1 \myifu/myicache/_2738_ ( .A(\myifu/myicache/_0647_ ), .B(\myifu/myicache/_0615_ ), .S(\myifu/myicache/_0949_ ), .Z(\myifu/myicache/_0338_ ) );
MUX2_X1 \myifu/myicache/_2739_ ( .A(\myifu/myicache/_0648_ ), .B(\myifu/myicache/_0616_ ), .S(\myifu/myicache/_0949_ ), .Z(\myifu/myicache/_0339_ ) );
AND2_X1 \myifu/myicache/_2740_ ( .A1(\myifu/myicache/_0900_ ), .A2(\myifu/myicache/_1228_ ), .ZN(\myifu/myicache/_0953_ ) );
MUX2_X1 \myifu/myicache/_2741_ ( .A(\myifu/myicache/_0953_ ), .B(\myifu/myicache/_1231_ ), .S(\myifu/myicache/_0945_ ), .Z(\myifu/myicache/_0340_ ) );
BUF_X4 \myifu/myicache/_2742_ ( .A(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0954_ ) );
MUX2_X1 \myifu/myicache/_2743_ ( .A(\myifu/myicache/_1146_ ), .B(\myifu/myicache/_1173_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0341_ ) );
MUX2_X1 \myifu/myicache/_2744_ ( .A(\myifu/myicache/_1157_ ), .B(\myifu/myicache/_1184_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0342_ ) );
MUX2_X1 \myifu/myicache/_2745_ ( .A(\myifu/myicache/_1165_ ), .B(\myifu/myicache/_1192_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0343_ ) );
MUX2_X1 \myifu/myicache/_2746_ ( .A(\myifu/myicache/_1166_ ), .B(\myifu/myicache/_1193_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0344_ ) );
MUX2_X1 \myifu/myicache/_2747_ ( .A(\myifu/myicache/_1167_ ), .B(\myifu/myicache/_1194_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0345_ ) );
MUX2_X1 \myifu/myicache/_2748_ ( .A(\myifu/myicache/_1168_ ), .B(\myifu/myicache/_1195_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0346_ ) );
MUX2_X1 \myifu/myicache/_2749_ ( .A(\myifu/myicache/_1169_ ), .B(\myifu/myicache/_1196_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0347_ ) );
MUX2_X1 \myifu/myicache/_2750_ ( .A(\myifu/myicache/_1170_ ), .B(\myifu/myicache/_1197_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0348_ ) );
MUX2_X1 \myifu/myicache/_2751_ ( .A(\myifu/myicache/_1171_ ), .B(\myifu/myicache/_1198_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0349_ ) );
MUX2_X1 \myifu/myicache/_2752_ ( .A(\myifu/myicache/_1172_ ), .B(\myifu/myicache/_1199_ ), .S(\myifu/myicache/_0954_ ), .Z(\myifu/myicache/_0350_ ) );
BUF_X4 \myifu/myicache/_2753_ ( .A(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0955_ ) );
MUX2_X1 \myifu/myicache/_2754_ ( .A(\myifu/myicache/_1147_ ), .B(\myifu/myicache/_1174_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0351_ ) );
MUX2_X1 \myifu/myicache/_2755_ ( .A(\myifu/myicache/_1148_ ), .B(\myifu/myicache/_1175_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0352_ ) );
MUX2_X1 \myifu/myicache/_2756_ ( .A(\myifu/myicache/_1149_ ), .B(\myifu/myicache/_1176_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0353_ ) );
MUX2_X1 \myifu/myicache/_2757_ ( .A(\myifu/myicache/_1150_ ), .B(\myifu/myicache/_1177_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0354_ ) );
MUX2_X1 \myifu/myicache/_2758_ ( .A(\myifu/myicache/_1151_ ), .B(\myifu/myicache/_1178_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0355_ ) );
MUX2_X1 \myifu/myicache/_2759_ ( .A(\myifu/myicache/_1152_ ), .B(\myifu/myicache/_1179_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0356_ ) );
MUX2_X1 \myifu/myicache/_2760_ ( .A(\myifu/myicache/_1153_ ), .B(\myifu/myicache/_1180_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0357_ ) );
MUX2_X1 \myifu/myicache/_2761_ ( .A(\myifu/myicache/_1154_ ), .B(\myifu/myicache/_1181_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0358_ ) );
MUX2_X1 \myifu/myicache/_2762_ ( .A(\myifu/myicache/_1155_ ), .B(\myifu/myicache/_1182_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0359_ ) );
MUX2_X1 \myifu/myicache/_2763_ ( .A(\myifu/myicache/_1156_ ), .B(\myifu/myicache/_1183_ ), .S(\myifu/myicache/_0955_ ), .Z(\myifu/myicache/_0360_ ) );
MUX2_X1 \myifu/myicache/_2764_ ( .A(\myifu/myicache/_1158_ ), .B(\myifu/myicache/_1185_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0361_ ) );
MUX2_X1 \myifu/myicache/_2765_ ( .A(\myifu/myicache/_1159_ ), .B(\myifu/myicache/_1186_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0362_ ) );
MUX2_X1 \myifu/myicache/_2766_ ( .A(\myifu/myicache/_1160_ ), .B(\myifu/myicache/_1187_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0363_ ) );
MUX2_X1 \myifu/myicache/_2767_ ( .A(\myifu/myicache/_1161_ ), .B(\myifu/myicache/_1188_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0364_ ) );
MUX2_X1 \myifu/myicache/_2768_ ( .A(\myifu/myicache/_1162_ ), .B(\myifu/myicache/_1189_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0365_ ) );
MUX2_X1 \myifu/myicache/_2769_ ( .A(\myifu/myicache/_1163_ ), .B(\myifu/myicache/_1190_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0366_ ) );
MUX2_X1 \myifu/myicache/_2770_ ( .A(\myifu/myicache/_1164_ ), .B(\myifu/myicache/_1191_ ), .S(\myifu/myicache/_0912_ ), .Z(\myifu/myicache/_0367_ ) );
DFF_X1 \myifu/myicache/_2771_ ( .D(\myifu/myicache/_1602_ ), .CK(clock ), .Q(\myifu/myicache/data[5][0] ), .QN(\myifu/myicache/_1601_ ) );
DFF_X1 \myifu/myicache/_2772_ ( .D(\myifu/myicache/_1603_ ), .CK(clock ), .Q(\myifu/myicache/data[5][1] ), .QN(\myifu/myicache/_1600_ ) );
DFF_X1 \myifu/myicache/_2773_ ( .D(\myifu/myicache/_1604_ ), .CK(clock ), .Q(\myifu/myicache/data[5][2] ), .QN(\myifu/myicache/_1599_ ) );
DFF_X1 \myifu/myicache/_2774_ ( .D(\myifu/myicache/_1605_ ), .CK(clock ), .Q(\myifu/myicache/data[5][3] ), .QN(\myifu/myicache/_1598_ ) );
DFF_X1 \myifu/myicache/_2775_ ( .D(\myifu/myicache/_1606_ ), .CK(clock ), .Q(\myifu/myicache/data[5][4] ), .QN(\myifu/myicache/_1597_ ) );
DFF_X1 \myifu/myicache/_2776_ ( .D(\myifu/myicache/_1607_ ), .CK(clock ), .Q(\myifu/myicache/data[5][5] ), .QN(\myifu/myicache/_1596_ ) );
DFF_X1 \myifu/myicache/_2777_ ( .D(\myifu/myicache/_1608_ ), .CK(clock ), .Q(\myifu/myicache/data[5][6] ), .QN(\myifu/myicache/_1595_ ) );
DFF_X1 \myifu/myicache/_2778_ ( .D(\myifu/myicache/_1609_ ), .CK(clock ), .Q(\myifu/myicache/data[5][7] ), .QN(\myifu/myicache/_1594_ ) );
DFF_X1 \myifu/myicache/_2779_ ( .D(\myifu/myicache/_1610_ ), .CK(clock ), .Q(\myifu/myicache/data[5][8] ), .QN(\myifu/myicache/_1593_ ) );
DFF_X1 \myifu/myicache/_2780_ ( .D(\myifu/myicache/_1611_ ), .CK(clock ), .Q(\myifu/myicache/data[5][9] ), .QN(\myifu/myicache/_1592_ ) );
DFF_X1 \myifu/myicache/_2781_ ( .D(\myifu/myicache/_1612_ ), .CK(clock ), .Q(\myifu/myicache/data[5][10] ), .QN(\myifu/myicache/_1591_ ) );
DFF_X1 \myifu/myicache/_2782_ ( .D(\myifu/myicache/_1613_ ), .CK(clock ), .Q(\myifu/myicache/data[5][11] ), .QN(\myifu/myicache/_1590_ ) );
DFF_X1 \myifu/myicache/_2783_ ( .D(\myifu/myicache/_1614_ ), .CK(clock ), .Q(\myifu/myicache/data[5][12] ), .QN(\myifu/myicache/_1589_ ) );
DFF_X1 \myifu/myicache/_2784_ ( .D(\myifu/myicache/_1615_ ), .CK(clock ), .Q(\myifu/myicache/data[5][13] ), .QN(\myifu/myicache/_1588_ ) );
DFF_X1 \myifu/myicache/_2785_ ( .D(\myifu/myicache/_1616_ ), .CK(clock ), .Q(\myifu/myicache/data[5][14] ), .QN(\myifu/myicache/_1587_ ) );
DFF_X1 \myifu/myicache/_2786_ ( .D(\myifu/myicache/_1617_ ), .CK(clock ), .Q(\myifu/myicache/data[5][15] ), .QN(\myifu/myicache/_1586_ ) );
DFF_X1 \myifu/myicache/_2787_ ( .D(\myifu/myicache/_1618_ ), .CK(clock ), .Q(\myifu/myicache/data[5][16] ), .QN(\myifu/myicache/_1585_ ) );
DFF_X1 \myifu/myicache/_2788_ ( .D(\myifu/myicache/_1619_ ), .CK(clock ), .Q(\myifu/myicache/data[5][17] ), .QN(\myifu/myicache/_1584_ ) );
DFF_X1 \myifu/myicache/_2789_ ( .D(\myifu/myicache/_1620_ ), .CK(clock ), .Q(\myifu/myicache/data[5][18] ), .QN(\myifu/myicache/_1583_ ) );
DFF_X1 \myifu/myicache/_2790_ ( .D(\myifu/myicache/_1621_ ), .CK(clock ), .Q(\myifu/myicache/data[5][19] ), .QN(\myifu/myicache/_1582_ ) );
DFF_X1 \myifu/myicache/_2791_ ( .D(\myifu/myicache/_1622_ ), .CK(clock ), .Q(\myifu/myicache/data[5][20] ), .QN(\myifu/myicache/_1581_ ) );
DFF_X1 \myifu/myicache/_2792_ ( .D(\myifu/myicache/_1623_ ), .CK(clock ), .Q(\myifu/myicache/data[5][21] ), .QN(\myifu/myicache/_1580_ ) );
DFF_X1 \myifu/myicache/_2793_ ( .D(\myifu/myicache/_1624_ ), .CK(clock ), .Q(\myifu/myicache/data[5][22] ), .QN(\myifu/myicache/_1579_ ) );
DFF_X1 \myifu/myicache/_2794_ ( .D(\myifu/myicache/_1625_ ), .CK(clock ), .Q(\myifu/myicache/data[5][23] ), .QN(\myifu/myicache/_1578_ ) );
DFF_X1 \myifu/myicache/_2795_ ( .D(\myifu/myicache/_1626_ ), .CK(clock ), .Q(\myifu/myicache/data[5][24] ), .QN(\myifu/myicache/_1577_ ) );
DFF_X1 \myifu/myicache/_2796_ ( .D(\myifu/myicache/_1627_ ), .CK(clock ), .Q(\myifu/myicache/data[5][25] ), .QN(\myifu/myicache/_1576_ ) );
DFF_X1 \myifu/myicache/_2797_ ( .D(\myifu/myicache/_1628_ ), .CK(clock ), .Q(\myifu/myicache/data[5][26] ), .QN(\myifu/myicache/_1575_ ) );
DFF_X1 \myifu/myicache/_2798_ ( .D(\myifu/myicache/_1629_ ), .CK(clock ), .Q(\myifu/myicache/data[5][27] ), .QN(\myifu/myicache/_1574_ ) );
DFF_X1 \myifu/myicache/_2799_ ( .D(\myifu/myicache/_1630_ ), .CK(clock ), .Q(\myifu/myicache/data[5][28] ), .QN(\myifu/myicache/_1573_ ) );
DFF_X1 \myifu/myicache/_2800_ ( .D(\myifu/myicache/_1631_ ), .CK(clock ), .Q(\myifu/myicache/data[5][29] ), .QN(\myifu/myicache/_1572_ ) );
DFF_X1 \myifu/myicache/_2801_ ( .D(\myifu/myicache/_1632_ ), .CK(clock ), .Q(\myifu/myicache/data[5][30] ), .QN(\myifu/myicache/_1571_ ) );
DFF_X1 \myifu/myicache/_2802_ ( .D(\myifu/myicache/_1633_ ), .CK(clock ), .Q(\myifu/myicache/data[5][31] ), .QN(\myifu/myicache/_1570_ ) );
DFF_X1 \myifu/myicache/_2803_ ( .D(\myifu/myicache/_1634_ ), .CK(clock ), .Q(\myifu/myicache/data[4][0] ), .QN(\myifu/myicache/_1569_ ) );
DFF_X1 \myifu/myicache/_2804_ ( .D(\myifu/myicache/_1635_ ), .CK(clock ), .Q(\myifu/myicache/data[4][1] ), .QN(\myifu/myicache/_1568_ ) );
DFF_X1 \myifu/myicache/_2805_ ( .D(\myifu/myicache/_1636_ ), .CK(clock ), .Q(\myifu/myicache/data[4][2] ), .QN(\myifu/myicache/_1567_ ) );
DFF_X1 \myifu/myicache/_2806_ ( .D(\myifu/myicache/_1637_ ), .CK(clock ), .Q(\myifu/myicache/data[4][3] ), .QN(\myifu/myicache/_1566_ ) );
DFF_X1 \myifu/myicache/_2807_ ( .D(\myifu/myicache/_1638_ ), .CK(clock ), .Q(\myifu/myicache/data[4][4] ), .QN(\myifu/myicache/_1565_ ) );
DFF_X1 \myifu/myicache/_2808_ ( .D(\myifu/myicache/_1639_ ), .CK(clock ), .Q(\myifu/myicache/data[4][5] ), .QN(\myifu/myicache/_1564_ ) );
DFF_X1 \myifu/myicache/_2809_ ( .D(\myifu/myicache/_1640_ ), .CK(clock ), .Q(\myifu/myicache/data[4][6] ), .QN(\myifu/myicache/_1563_ ) );
DFF_X1 \myifu/myicache/_2810_ ( .D(\myifu/myicache/_1641_ ), .CK(clock ), .Q(\myifu/myicache/data[4][7] ), .QN(\myifu/myicache/_1562_ ) );
DFF_X1 \myifu/myicache/_2811_ ( .D(\myifu/myicache/_1642_ ), .CK(clock ), .Q(\myifu/myicache/data[4][8] ), .QN(\myifu/myicache/_1561_ ) );
DFF_X1 \myifu/myicache/_2812_ ( .D(\myifu/myicache/_1643_ ), .CK(clock ), .Q(\myifu/myicache/data[4][9] ), .QN(\myifu/myicache/_1560_ ) );
DFF_X1 \myifu/myicache/_2813_ ( .D(\myifu/myicache/_1644_ ), .CK(clock ), .Q(\myifu/myicache/data[4][10] ), .QN(\myifu/myicache/_1559_ ) );
DFF_X1 \myifu/myicache/_2814_ ( .D(\myifu/myicache/_1645_ ), .CK(clock ), .Q(\myifu/myicache/data[4][11] ), .QN(\myifu/myicache/_1558_ ) );
DFF_X1 \myifu/myicache/_2815_ ( .D(\myifu/myicache/_1646_ ), .CK(clock ), .Q(\myifu/myicache/data[4][12] ), .QN(\myifu/myicache/_1557_ ) );
DFF_X1 \myifu/myicache/_2816_ ( .D(\myifu/myicache/_1647_ ), .CK(clock ), .Q(\myifu/myicache/data[4][13] ), .QN(\myifu/myicache/_1556_ ) );
DFF_X1 \myifu/myicache/_2817_ ( .D(\myifu/myicache/_1648_ ), .CK(clock ), .Q(\myifu/myicache/data[4][14] ), .QN(\myifu/myicache/_1555_ ) );
DFF_X1 \myifu/myicache/_2818_ ( .D(\myifu/myicache/_1649_ ), .CK(clock ), .Q(\myifu/myicache/data[4][15] ), .QN(\myifu/myicache/_1554_ ) );
DFF_X1 \myifu/myicache/_2819_ ( .D(\myifu/myicache/_1650_ ), .CK(clock ), .Q(\myifu/myicache/data[4][16] ), .QN(\myifu/myicache/_1553_ ) );
DFF_X1 \myifu/myicache/_2820_ ( .D(\myifu/myicache/_1651_ ), .CK(clock ), .Q(\myifu/myicache/data[4][17] ), .QN(\myifu/myicache/_1552_ ) );
DFF_X1 \myifu/myicache/_2821_ ( .D(\myifu/myicache/_1652_ ), .CK(clock ), .Q(\myifu/myicache/data[4][18] ), .QN(\myifu/myicache/_1551_ ) );
DFF_X1 \myifu/myicache/_2822_ ( .D(\myifu/myicache/_1653_ ), .CK(clock ), .Q(\myifu/myicache/data[4][19] ), .QN(\myifu/myicache/_1550_ ) );
DFF_X1 \myifu/myicache/_2823_ ( .D(\myifu/myicache/_1654_ ), .CK(clock ), .Q(\myifu/myicache/data[4][20] ), .QN(\myifu/myicache/_1549_ ) );
DFF_X1 \myifu/myicache/_2824_ ( .D(\myifu/myicache/_1655_ ), .CK(clock ), .Q(\myifu/myicache/data[4][21] ), .QN(\myifu/myicache/_1548_ ) );
DFF_X1 \myifu/myicache/_2825_ ( .D(\myifu/myicache/_1656_ ), .CK(clock ), .Q(\myifu/myicache/data[4][22] ), .QN(\myifu/myicache/_1547_ ) );
DFF_X1 \myifu/myicache/_2826_ ( .D(\myifu/myicache/_1657_ ), .CK(clock ), .Q(\myifu/myicache/data[4][23] ), .QN(\myifu/myicache/_1546_ ) );
DFF_X1 \myifu/myicache/_2827_ ( .D(\myifu/myicache/_1658_ ), .CK(clock ), .Q(\myifu/myicache/data[4][24] ), .QN(\myifu/myicache/_1545_ ) );
DFF_X1 \myifu/myicache/_2828_ ( .D(\myifu/myicache/_1659_ ), .CK(clock ), .Q(\myifu/myicache/data[4][25] ), .QN(\myifu/myicache/_1544_ ) );
DFF_X1 \myifu/myicache/_2829_ ( .D(\myifu/myicache/_1660_ ), .CK(clock ), .Q(\myifu/myicache/data[4][26] ), .QN(\myifu/myicache/_1543_ ) );
DFF_X1 \myifu/myicache/_2830_ ( .D(\myifu/myicache/_1661_ ), .CK(clock ), .Q(\myifu/myicache/data[4][27] ), .QN(\myifu/myicache/_1542_ ) );
DFF_X1 \myifu/myicache/_2831_ ( .D(\myifu/myicache/_1662_ ), .CK(clock ), .Q(\myifu/myicache/data[4][28] ), .QN(\myifu/myicache/_1541_ ) );
DFF_X1 \myifu/myicache/_2832_ ( .D(\myifu/myicache/_1663_ ), .CK(clock ), .Q(\myifu/myicache/data[4][29] ), .QN(\myifu/myicache/_1540_ ) );
DFF_X1 \myifu/myicache/_2833_ ( .D(\myifu/myicache/_1664_ ), .CK(clock ), .Q(\myifu/myicache/data[4][30] ), .QN(\myifu/myicache/_1539_ ) );
DFF_X1 \myifu/myicache/_2834_ ( .D(\myifu/myicache/_1665_ ), .CK(clock ), .Q(\myifu/myicache/data[4][31] ), .QN(\myifu/myicache/_1538_ ) );
DFF_X1 \myifu/myicache/_2835_ ( .D(\myifu/myicache/_1666_ ), .CK(clock ), .Q(\myifu/myicache/data[6][0] ), .QN(\myifu/myicache/_1537_ ) );
DFF_X1 \myifu/myicache/_2836_ ( .D(\myifu/myicache/_1667_ ), .CK(clock ), .Q(\myifu/myicache/data[6][1] ), .QN(\myifu/myicache/_1536_ ) );
DFF_X1 \myifu/myicache/_2837_ ( .D(\myifu/myicache/_1668_ ), .CK(clock ), .Q(\myifu/myicache/data[6][2] ), .QN(\myifu/myicache/_1535_ ) );
DFF_X1 \myifu/myicache/_2838_ ( .D(\myifu/myicache/_1669_ ), .CK(clock ), .Q(\myifu/myicache/data[6][3] ), .QN(\myifu/myicache/_1534_ ) );
DFF_X1 \myifu/myicache/_2839_ ( .D(\myifu/myicache/_1670_ ), .CK(clock ), .Q(\myifu/myicache/data[6][4] ), .QN(\myifu/myicache/_1533_ ) );
DFF_X1 \myifu/myicache/_2840_ ( .D(\myifu/myicache/_1671_ ), .CK(clock ), .Q(\myifu/myicache/data[6][5] ), .QN(\myifu/myicache/_1532_ ) );
DFF_X1 \myifu/myicache/_2841_ ( .D(\myifu/myicache/_1672_ ), .CK(clock ), .Q(\myifu/myicache/data[6][6] ), .QN(\myifu/myicache/_1531_ ) );
DFF_X1 \myifu/myicache/_2842_ ( .D(\myifu/myicache/_1673_ ), .CK(clock ), .Q(\myifu/myicache/data[6][7] ), .QN(\myifu/myicache/_1530_ ) );
DFF_X1 \myifu/myicache/_2843_ ( .D(\myifu/myicache/_1674_ ), .CK(clock ), .Q(\myifu/myicache/data[6][8] ), .QN(\myifu/myicache/_1529_ ) );
DFF_X1 \myifu/myicache/_2844_ ( .D(\myifu/myicache/_1675_ ), .CK(clock ), .Q(\myifu/myicache/data[6][9] ), .QN(\myifu/myicache/_1528_ ) );
DFF_X1 \myifu/myicache/_2845_ ( .D(\myifu/myicache/_1676_ ), .CK(clock ), .Q(\myifu/myicache/data[6][10] ), .QN(\myifu/myicache/_1527_ ) );
DFF_X1 \myifu/myicache/_2846_ ( .D(\myifu/myicache/_1677_ ), .CK(clock ), .Q(\myifu/myicache/data[6][11] ), .QN(\myifu/myicache/_1526_ ) );
DFF_X1 \myifu/myicache/_2847_ ( .D(\myifu/myicache/_1678_ ), .CK(clock ), .Q(\myifu/myicache/data[6][12] ), .QN(\myifu/myicache/_1525_ ) );
DFF_X1 \myifu/myicache/_2848_ ( .D(\myifu/myicache/_1679_ ), .CK(clock ), .Q(\myifu/myicache/data[6][13] ), .QN(\myifu/myicache/_1524_ ) );
DFF_X1 \myifu/myicache/_2849_ ( .D(\myifu/myicache/_1680_ ), .CK(clock ), .Q(\myifu/myicache/data[6][14] ), .QN(\myifu/myicache/_1523_ ) );
DFF_X1 \myifu/myicache/_2850_ ( .D(\myifu/myicache/_1681_ ), .CK(clock ), .Q(\myifu/myicache/data[6][15] ), .QN(\myifu/myicache/_1522_ ) );
DFF_X1 \myifu/myicache/_2851_ ( .D(\myifu/myicache/_1682_ ), .CK(clock ), .Q(\myifu/myicache/data[6][16] ), .QN(\myifu/myicache/_1521_ ) );
DFF_X1 \myifu/myicache/_2852_ ( .D(\myifu/myicache/_1683_ ), .CK(clock ), .Q(\myifu/myicache/data[6][17] ), .QN(\myifu/myicache/_1520_ ) );
DFF_X1 \myifu/myicache/_2853_ ( .D(\myifu/myicache/_1684_ ), .CK(clock ), .Q(\myifu/myicache/data[6][18] ), .QN(\myifu/myicache/_1519_ ) );
DFF_X1 \myifu/myicache/_2854_ ( .D(\myifu/myicache/_1685_ ), .CK(clock ), .Q(\myifu/myicache/data[6][19] ), .QN(\myifu/myicache/_1518_ ) );
DFF_X1 \myifu/myicache/_2855_ ( .D(\myifu/myicache/_1686_ ), .CK(clock ), .Q(\myifu/myicache/data[6][20] ), .QN(\myifu/myicache/_1517_ ) );
DFF_X1 \myifu/myicache/_2856_ ( .D(\myifu/myicache/_1687_ ), .CK(clock ), .Q(\myifu/myicache/data[6][21] ), .QN(\myifu/myicache/_1516_ ) );
DFF_X1 \myifu/myicache/_2857_ ( .D(\myifu/myicache/_1688_ ), .CK(clock ), .Q(\myifu/myicache/data[6][22] ), .QN(\myifu/myicache/_1515_ ) );
DFF_X1 \myifu/myicache/_2858_ ( .D(\myifu/myicache/_1689_ ), .CK(clock ), .Q(\myifu/myicache/data[6][23] ), .QN(\myifu/myicache/_1514_ ) );
DFF_X1 \myifu/myicache/_2859_ ( .D(\myifu/myicache/_1690_ ), .CK(clock ), .Q(\myifu/myicache/data[6][24] ), .QN(\myifu/myicache/_1513_ ) );
DFF_X1 \myifu/myicache/_2860_ ( .D(\myifu/myicache/_1691_ ), .CK(clock ), .Q(\myifu/myicache/data[6][25] ), .QN(\myifu/myicache/_1512_ ) );
DFF_X1 \myifu/myicache/_2861_ ( .D(\myifu/myicache/_1692_ ), .CK(clock ), .Q(\myifu/myicache/data[6][26] ), .QN(\myifu/myicache/_1511_ ) );
DFF_X1 \myifu/myicache/_2862_ ( .D(\myifu/myicache/_1693_ ), .CK(clock ), .Q(\myifu/myicache/data[6][27] ), .QN(\myifu/myicache/_1510_ ) );
DFF_X1 \myifu/myicache/_2863_ ( .D(\myifu/myicache/_1694_ ), .CK(clock ), .Q(\myifu/myicache/data[6][28] ), .QN(\myifu/myicache/_1509_ ) );
DFF_X1 \myifu/myicache/_2864_ ( .D(\myifu/myicache/_1695_ ), .CK(clock ), .Q(\myifu/myicache/data[6][29] ), .QN(\myifu/myicache/_1508_ ) );
DFF_X1 \myifu/myicache/_2865_ ( .D(\myifu/myicache/_1696_ ), .CK(clock ), .Q(\myifu/myicache/data[6][30] ), .QN(\myifu/myicache/_1507_ ) );
DFF_X1 \myifu/myicache/_2866_ ( .D(\myifu/myicache/_1697_ ), .CK(clock ), .Q(\myifu/myicache/data[6][31] ), .QN(\myifu/myicache/_1506_ ) );
DFF_X1 \myifu/myicache/_2867_ ( .D(\myifu/myicache/_1698_ ), .CK(clock ), .Q(\myifu/myicache/valid [2] ), .QN(\myifu/myicache/_1505_ ) );
DFF_X1 \myifu/myicache/_2868_ ( .D(\myifu/myicache/_1699_ ), .CK(clock ), .Q(\myifu/myicache/valid [0] ), .QN(\myifu/myicache/_1504_ ) );
DFF_X1 \myifu/myicache/_2869_ ( .D(\myifu/myicache/_1700_ ), .CK(clock ), .Q(\myifu/myicache/data[2][0] ), .QN(\myifu/myicache/_1503_ ) );
DFF_X1 \myifu/myicache/_2870_ ( .D(\myifu/myicache/_1701_ ), .CK(clock ), .Q(\myifu/myicache/data[2][1] ), .QN(\myifu/myicache/_1502_ ) );
DFF_X1 \myifu/myicache/_2871_ ( .D(\myifu/myicache/_1702_ ), .CK(clock ), .Q(\myifu/myicache/data[2][2] ), .QN(\myifu/myicache/_1501_ ) );
DFF_X1 \myifu/myicache/_2872_ ( .D(\myifu/myicache/_1703_ ), .CK(clock ), .Q(\myifu/myicache/data[2][3] ), .QN(\myifu/myicache/_1500_ ) );
DFF_X1 \myifu/myicache/_2873_ ( .D(\myifu/myicache/_1704_ ), .CK(clock ), .Q(\myifu/myicache/data[2][4] ), .QN(\myifu/myicache/_1499_ ) );
DFF_X1 \myifu/myicache/_2874_ ( .D(\myifu/myicache/_1705_ ), .CK(clock ), .Q(\myifu/myicache/data[2][5] ), .QN(\myifu/myicache/_1498_ ) );
DFF_X1 \myifu/myicache/_2875_ ( .D(\myifu/myicache/_1706_ ), .CK(clock ), .Q(\myifu/myicache/data[2][6] ), .QN(\myifu/myicache/_1497_ ) );
DFF_X1 \myifu/myicache/_2876_ ( .D(\myifu/myicache/_1707_ ), .CK(clock ), .Q(\myifu/myicache/data[2][7] ), .QN(\myifu/myicache/_1496_ ) );
DFF_X1 \myifu/myicache/_2877_ ( .D(\myifu/myicache/_1708_ ), .CK(clock ), .Q(\myifu/myicache/data[2][8] ), .QN(\myifu/myicache/_1495_ ) );
DFF_X1 \myifu/myicache/_2878_ ( .D(\myifu/myicache/_1709_ ), .CK(clock ), .Q(\myifu/myicache/data[2][9] ), .QN(\myifu/myicache/_1494_ ) );
DFF_X1 \myifu/myicache/_2879_ ( .D(\myifu/myicache/_1710_ ), .CK(clock ), .Q(\myifu/myicache/data[2][10] ), .QN(\myifu/myicache/_1493_ ) );
DFF_X1 \myifu/myicache/_2880_ ( .D(\myifu/myicache/_1711_ ), .CK(clock ), .Q(\myifu/myicache/data[2][11] ), .QN(\myifu/myicache/_1492_ ) );
DFF_X1 \myifu/myicache/_2881_ ( .D(\myifu/myicache/_1712_ ), .CK(clock ), .Q(\myifu/myicache/data[2][12] ), .QN(\myifu/myicache/_1491_ ) );
DFF_X1 \myifu/myicache/_2882_ ( .D(\myifu/myicache/_1713_ ), .CK(clock ), .Q(\myifu/myicache/data[2][13] ), .QN(\myifu/myicache/_1490_ ) );
DFF_X1 \myifu/myicache/_2883_ ( .D(\myifu/myicache/_1714_ ), .CK(clock ), .Q(\myifu/myicache/data[2][14] ), .QN(\myifu/myicache/_1489_ ) );
DFF_X1 \myifu/myicache/_2884_ ( .D(\myifu/myicache/_1715_ ), .CK(clock ), .Q(\myifu/myicache/data[2][15] ), .QN(\myifu/myicache/_1488_ ) );
DFF_X1 \myifu/myicache/_2885_ ( .D(\myifu/myicache/_1716_ ), .CK(clock ), .Q(\myifu/myicache/data[2][16] ), .QN(\myifu/myicache/_1487_ ) );
DFF_X1 \myifu/myicache/_2886_ ( .D(\myifu/myicache/_1717_ ), .CK(clock ), .Q(\myifu/myicache/data[2][17] ), .QN(\myifu/myicache/_1486_ ) );
DFF_X1 \myifu/myicache/_2887_ ( .D(\myifu/myicache/_1718_ ), .CK(clock ), .Q(\myifu/myicache/data[2][18] ), .QN(\myifu/myicache/_1485_ ) );
DFF_X1 \myifu/myicache/_2888_ ( .D(\myifu/myicache/_1719_ ), .CK(clock ), .Q(\myifu/myicache/data[2][19] ), .QN(\myifu/myicache/_1484_ ) );
DFF_X1 \myifu/myicache/_2889_ ( .D(\myifu/myicache/_1720_ ), .CK(clock ), .Q(\myifu/myicache/data[2][20] ), .QN(\myifu/myicache/_1483_ ) );
DFF_X1 \myifu/myicache/_2890_ ( .D(\myifu/myicache/_1721_ ), .CK(clock ), .Q(\myifu/myicache/data[2][21] ), .QN(\myifu/myicache/_1482_ ) );
DFF_X1 \myifu/myicache/_2891_ ( .D(\myifu/myicache/_1722_ ), .CK(clock ), .Q(\myifu/myicache/data[2][22] ), .QN(\myifu/myicache/_1481_ ) );
DFF_X1 \myifu/myicache/_2892_ ( .D(\myifu/myicache/_1723_ ), .CK(clock ), .Q(\myifu/myicache/data[2][23] ), .QN(\myifu/myicache/_1480_ ) );
DFF_X1 \myifu/myicache/_2893_ ( .D(\myifu/myicache/_1724_ ), .CK(clock ), .Q(\myifu/myicache/data[2][24] ), .QN(\myifu/myicache/_1479_ ) );
DFF_X1 \myifu/myicache/_2894_ ( .D(\myifu/myicache/_1725_ ), .CK(clock ), .Q(\myifu/myicache/data[2][25] ), .QN(\myifu/myicache/_1478_ ) );
DFF_X1 \myifu/myicache/_2895_ ( .D(\myifu/myicache/_1726_ ), .CK(clock ), .Q(\myifu/myicache/data[2][26] ), .QN(\myifu/myicache/_1477_ ) );
DFF_X1 \myifu/myicache/_2896_ ( .D(\myifu/myicache/_1727_ ), .CK(clock ), .Q(\myifu/myicache/data[2][27] ), .QN(\myifu/myicache/_1476_ ) );
DFF_X1 \myifu/myicache/_2897_ ( .D(\myifu/myicache/_1728_ ), .CK(clock ), .Q(\myifu/myicache/data[2][28] ), .QN(\myifu/myicache/_1475_ ) );
DFF_X1 \myifu/myicache/_2898_ ( .D(\myifu/myicache/_1729_ ), .CK(clock ), .Q(\myifu/myicache/data[2][29] ), .QN(\myifu/myicache/_1474_ ) );
DFF_X1 \myifu/myicache/_2899_ ( .D(\myifu/myicache/_1730_ ), .CK(clock ), .Q(\myifu/myicache/data[2][30] ), .QN(\myifu/myicache/_1473_ ) );
DFF_X1 \myifu/myicache/_2900_ ( .D(\myifu/myicache/_1731_ ), .CK(clock ), .Q(\myifu/myicache/data[2][31] ), .QN(\myifu/myicache/_1472_ ) );
DFF_X1 \myifu/myicache/_2901_ ( .D(\myifu/myicache/_1732_ ), .CK(clock ), .Q(\myifu/myicache/data[1][0] ), .QN(\myifu/myicache/_1471_ ) );
DFF_X1 \myifu/myicache/_2902_ ( .D(\myifu/myicache/_1733_ ), .CK(clock ), .Q(\myifu/myicache/data[1][1] ), .QN(\myifu/myicache/_1470_ ) );
DFF_X1 \myifu/myicache/_2903_ ( .D(\myifu/myicache/_1734_ ), .CK(clock ), .Q(\myifu/myicache/data[1][2] ), .QN(\myifu/myicache/_1469_ ) );
DFF_X1 \myifu/myicache/_2904_ ( .D(\myifu/myicache/_1735_ ), .CK(clock ), .Q(\myifu/myicache/data[1][3] ), .QN(\myifu/myicache/_1468_ ) );
DFF_X1 \myifu/myicache/_2905_ ( .D(\myifu/myicache/_1736_ ), .CK(clock ), .Q(\myifu/myicache/data[1][4] ), .QN(\myifu/myicache/_1467_ ) );
DFF_X1 \myifu/myicache/_2906_ ( .D(\myifu/myicache/_1737_ ), .CK(clock ), .Q(\myifu/myicache/data[1][5] ), .QN(\myifu/myicache/_1466_ ) );
DFF_X1 \myifu/myicache/_2907_ ( .D(\myifu/myicache/_1738_ ), .CK(clock ), .Q(\myifu/myicache/data[1][6] ), .QN(\myifu/myicache/_1465_ ) );
DFF_X1 \myifu/myicache/_2908_ ( .D(\myifu/myicache/_1739_ ), .CK(clock ), .Q(\myifu/myicache/data[1][7] ), .QN(\myifu/myicache/_1464_ ) );
DFF_X1 \myifu/myicache/_2909_ ( .D(\myifu/myicache/_1740_ ), .CK(clock ), .Q(\myifu/myicache/data[1][8] ), .QN(\myifu/myicache/_1463_ ) );
DFF_X1 \myifu/myicache/_2910_ ( .D(\myifu/myicache/_1741_ ), .CK(clock ), .Q(\myifu/myicache/data[1][9] ), .QN(\myifu/myicache/_1462_ ) );
DFF_X1 \myifu/myicache/_2911_ ( .D(\myifu/myicache/_1742_ ), .CK(clock ), .Q(\myifu/myicache/data[1][10] ), .QN(\myifu/myicache/_1461_ ) );
DFF_X1 \myifu/myicache/_2912_ ( .D(\myifu/myicache/_1743_ ), .CK(clock ), .Q(\myifu/myicache/data[1][11] ), .QN(\myifu/myicache/_1460_ ) );
DFF_X1 \myifu/myicache/_2913_ ( .D(\myifu/myicache/_1744_ ), .CK(clock ), .Q(\myifu/myicache/data[1][12] ), .QN(\myifu/myicache/_1459_ ) );
DFF_X1 \myifu/myicache/_2914_ ( .D(\myifu/myicache/_1745_ ), .CK(clock ), .Q(\myifu/myicache/data[1][13] ), .QN(\myifu/myicache/_1458_ ) );
DFF_X1 \myifu/myicache/_2915_ ( .D(\myifu/myicache/_1746_ ), .CK(clock ), .Q(\myifu/myicache/data[1][14] ), .QN(\myifu/myicache/_1457_ ) );
DFF_X1 \myifu/myicache/_2916_ ( .D(\myifu/myicache/_1747_ ), .CK(clock ), .Q(\myifu/myicache/data[1][15] ), .QN(\myifu/myicache/_1456_ ) );
DFF_X1 \myifu/myicache/_2917_ ( .D(\myifu/myicache/_1748_ ), .CK(clock ), .Q(\myifu/myicache/data[1][16] ), .QN(\myifu/myicache/_1455_ ) );
DFF_X1 \myifu/myicache/_2918_ ( .D(\myifu/myicache/_1749_ ), .CK(clock ), .Q(\myifu/myicache/data[1][17] ), .QN(\myifu/myicache/_1454_ ) );
DFF_X1 \myifu/myicache/_2919_ ( .D(\myifu/myicache/_1750_ ), .CK(clock ), .Q(\myifu/myicache/data[1][18] ), .QN(\myifu/myicache/_1453_ ) );
DFF_X1 \myifu/myicache/_2920_ ( .D(\myifu/myicache/_1751_ ), .CK(clock ), .Q(\myifu/myicache/data[1][19] ), .QN(\myifu/myicache/_1452_ ) );
DFF_X1 \myifu/myicache/_2921_ ( .D(\myifu/myicache/_1752_ ), .CK(clock ), .Q(\myifu/myicache/data[1][20] ), .QN(\myifu/myicache/_1451_ ) );
DFF_X1 \myifu/myicache/_2922_ ( .D(\myifu/myicache/_1753_ ), .CK(clock ), .Q(\myifu/myicache/data[1][21] ), .QN(\myifu/myicache/_1450_ ) );
DFF_X1 \myifu/myicache/_2923_ ( .D(\myifu/myicache/_1754_ ), .CK(clock ), .Q(\myifu/myicache/data[1][22] ), .QN(\myifu/myicache/_1449_ ) );
DFF_X1 \myifu/myicache/_2924_ ( .D(\myifu/myicache/_1755_ ), .CK(clock ), .Q(\myifu/myicache/data[1][23] ), .QN(\myifu/myicache/_1448_ ) );
DFF_X1 \myifu/myicache/_2925_ ( .D(\myifu/myicache/_1756_ ), .CK(clock ), .Q(\myifu/myicache/data[1][24] ), .QN(\myifu/myicache/_1447_ ) );
DFF_X1 \myifu/myicache/_2926_ ( .D(\myifu/myicache/_1757_ ), .CK(clock ), .Q(\myifu/myicache/data[1][25] ), .QN(\myifu/myicache/_1446_ ) );
DFF_X1 \myifu/myicache/_2927_ ( .D(\myifu/myicache/_1758_ ), .CK(clock ), .Q(\myifu/myicache/data[1][26] ), .QN(\myifu/myicache/_1445_ ) );
DFF_X1 \myifu/myicache/_2928_ ( .D(\myifu/myicache/_1759_ ), .CK(clock ), .Q(\myifu/myicache/data[1][27] ), .QN(\myifu/myicache/_1444_ ) );
DFF_X1 \myifu/myicache/_2929_ ( .D(\myifu/myicache/_1760_ ), .CK(clock ), .Q(\myifu/myicache/data[1][28] ), .QN(\myifu/myicache/_1443_ ) );
DFF_X1 \myifu/myicache/_2930_ ( .D(\myifu/myicache/_1761_ ), .CK(clock ), .Q(\myifu/myicache/data[1][29] ), .QN(\myifu/myicache/_1442_ ) );
DFF_X1 \myifu/myicache/_2931_ ( .D(\myifu/myicache/_1762_ ), .CK(clock ), .Q(\myifu/myicache/data[1][30] ), .QN(\myifu/myicache/_1441_ ) );
DFF_X1 \myifu/myicache/_2932_ ( .D(\myifu/myicache/_1763_ ), .CK(clock ), .Q(\myifu/myicache/data[1][31] ), .QN(\myifu/myicache/_1440_ ) );
DFF_X1 \myifu/myicache/_2933_ ( .D(\myifu/myicache/_1764_ ), .CK(clock ), .Q(\myifu/myicache/data[0][0] ), .QN(\myifu/myicache/_1439_ ) );
DFF_X1 \myifu/myicache/_2934_ ( .D(\myifu/myicache/_1765_ ), .CK(clock ), .Q(\myifu/myicache/data[0][1] ), .QN(\myifu/myicache/_1438_ ) );
DFF_X1 \myifu/myicache/_2935_ ( .D(\myifu/myicache/_1766_ ), .CK(clock ), .Q(\myifu/myicache/data[0][2] ), .QN(\myifu/myicache/_1437_ ) );
DFF_X1 \myifu/myicache/_2936_ ( .D(\myifu/myicache/_1767_ ), .CK(clock ), .Q(\myifu/myicache/data[0][3] ), .QN(\myifu/myicache/_1436_ ) );
DFF_X1 \myifu/myicache/_2937_ ( .D(\myifu/myicache/_1768_ ), .CK(clock ), .Q(\myifu/myicache/data[0][4] ), .QN(\myifu/myicache/_1435_ ) );
DFF_X1 \myifu/myicache/_2938_ ( .D(\myifu/myicache/_1769_ ), .CK(clock ), .Q(\myifu/myicache/data[0][5] ), .QN(\myifu/myicache/_1434_ ) );
DFF_X1 \myifu/myicache/_2939_ ( .D(\myifu/myicache/_1770_ ), .CK(clock ), .Q(\myifu/myicache/data[0][6] ), .QN(\myifu/myicache/_1433_ ) );
DFF_X1 \myifu/myicache/_2940_ ( .D(\myifu/myicache/_1771_ ), .CK(clock ), .Q(\myifu/myicache/data[0][7] ), .QN(\myifu/myicache/_1432_ ) );
DFF_X1 \myifu/myicache/_2941_ ( .D(\myifu/myicache/_1772_ ), .CK(clock ), .Q(\myifu/myicache/data[0][8] ), .QN(\myifu/myicache/_1431_ ) );
DFF_X1 \myifu/myicache/_2942_ ( .D(\myifu/myicache/_1773_ ), .CK(clock ), .Q(\myifu/myicache/data[0][9] ), .QN(\myifu/myicache/_1430_ ) );
DFF_X1 \myifu/myicache/_2943_ ( .D(\myifu/myicache/_1774_ ), .CK(clock ), .Q(\myifu/myicache/data[0][10] ), .QN(\myifu/myicache/_1429_ ) );
DFF_X1 \myifu/myicache/_2944_ ( .D(\myifu/myicache/_1775_ ), .CK(clock ), .Q(\myifu/myicache/data[0][11] ), .QN(\myifu/myicache/_1428_ ) );
DFF_X1 \myifu/myicache/_2945_ ( .D(\myifu/myicache/_1776_ ), .CK(clock ), .Q(\myifu/myicache/data[0][12] ), .QN(\myifu/myicache/_1427_ ) );
DFF_X1 \myifu/myicache/_2946_ ( .D(\myifu/myicache/_1777_ ), .CK(clock ), .Q(\myifu/myicache/data[0][13] ), .QN(\myifu/myicache/_1426_ ) );
DFF_X1 \myifu/myicache/_2947_ ( .D(\myifu/myicache/_1778_ ), .CK(clock ), .Q(\myifu/myicache/data[0][14] ), .QN(\myifu/myicache/_1425_ ) );
DFF_X1 \myifu/myicache/_2948_ ( .D(\myifu/myicache/_1779_ ), .CK(clock ), .Q(\myifu/myicache/data[0][15] ), .QN(\myifu/myicache/_1424_ ) );
DFF_X1 \myifu/myicache/_2949_ ( .D(\myifu/myicache/_1780_ ), .CK(clock ), .Q(\myifu/myicache/data[0][16] ), .QN(\myifu/myicache/_1423_ ) );
DFF_X1 \myifu/myicache/_2950_ ( .D(\myifu/myicache/_1781_ ), .CK(clock ), .Q(\myifu/myicache/data[0][17] ), .QN(\myifu/myicache/_1422_ ) );
DFF_X1 \myifu/myicache/_2951_ ( .D(\myifu/myicache/_1782_ ), .CK(clock ), .Q(\myifu/myicache/data[0][18] ), .QN(\myifu/myicache/_1421_ ) );
DFF_X1 \myifu/myicache/_2952_ ( .D(\myifu/myicache/_1783_ ), .CK(clock ), .Q(\myifu/myicache/data[0][19] ), .QN(\myifu/myicache/_1420_ ) );
DFF_X1 \myifu/myicache/_2953_ ( .D(\myifu/myicache/_1784_ ), .CK(clock ), .Q(\myifu/myicache/data[0][20] ), .QN(\myifu/myicache/_1419_ ) );
DFF_X1 \myifu/myicache/_2954_ ( .D(\myifu/myicache/_1785_ ), .CK(clock ), .Q(\myifu/myicache/data[0][21] ), .QN(\myifu/myicache/_1418_ ) );
DFF_X1 \myifu/myicache/_2955_ ( .D(\myifu/myicache/_1786_ ), .CK(clock ), .Q(\myifu/myicache/data[0][22] ), .QN(\myifu/myicache/_1417_ ) );
DFF_X1 \myifu/myicache/_2956_ ( .D(\myifu/myicache/_1787_ ), .CK(clock ), .Q(\myifu/myicache/data[0][23] ), .QN(\myifu/myicache/_1416_ ) );
DFF_X1 \myifu/myicache/_2957_ ( .D(\myifu/myicache/_1788_ ), .CK(clock ), .Q(\myifu/myicache/data[0][24] ), .QN(\myifu/myicache/_1415_ ) );
DFF_X1 \myifu/myicache/_2958_ ( .D(\myifu/myicache/_1789_ ), .CK(clock ), .Q(\myifu/myicache/data[0][25] ), .QN(\myifu/myicache/_1414_ ) );
DFF_X1 \myifu/myicache/_2959_ ( .D(\myifu/myicache/_1790_ ), .CK(clock ), .Q(\myifu/myicache/data[0][26] ), .QN(\myifu/myicache/_1413_ ) );
DFF_X1 \myifu/myicache/_2960_ ( .D(\myifu/myicache/_1791_ ), .CK(clock ), .Q(\myifu/myicache/data[0][27] ), .QN(\myifu/myicache/_1412_ ) );
DFF_X1 \myifu/myicache/_2961_ ( .D(\myifu/myicache/_1792_ ), .CK(clock ), .Q(\myifu/myicache/data[0][28] ), .QN(\myifu/myicache/_1411_ ) );
DFF_X1 \myifu/myicache/_2962_ ( .D(\myifu/myicache/_1793_ ), .CK(clock ), .Q(\myifu/myicache/data[0][29] ), .QN(\myifu/myicache/_1410_ ) );
DFF_X1 \myifu/myicache/_2963_ ( .D(\myifu/myicache/_1794_ ), .CK(clock ), .Q(\myifu/myicache/data[0][30] ), .QN(\myifu/myicache/_1409_ ) );
DFF_X1 \myifu/myicache/_2964_ ( .D(\myifu/myicache/_1795_ ), .CK(clock ), .Q(\myifu/myicache/data[0][31] ), .QN(\myifu/myicache/_1408_ ) );
DFF_X1 \myifu/myicache/_2965_ ( .D(\myifu/myicache/_1796_ ), .CK(clock ), .Q(\myifu/myicache/valid [3] ), .QN(\myifu/myicache/_1407_ ) );
DFF_X1 \myifu/myicache/_2966_ ( .D(\myifu/myicache/_1797_ ), .CK(clock ), .Q(\myifu/myicache/data[3][0] ), .QN(\myifu/myicache/_1406_ ) );
DFF_X1 \myifu/myicache/_2967_ ( .D(\myifu/myicache/_1798_ ), .CK(clock ), .Q(\myifu/myicache/data[3][1] ), .QN(\myifu/myicache/_1405_ ) );
DFF_X1 \myifu/myicache/_2968_ ( .D(\myifu/myicache/_1799_ ), .CK(clock ), .Q(\myifu/myicache/data[3][2] ), .QN(\myifu/myicache/_1404_ ) );
DFF_X1 \myifu/myicache/_2969_ ( .D(\myifu/myicache/_1800_ ), .CK(clock ), .Q(\myifu/myicache/data[3][3] ), .QN(\myifu/myicache/_1403_ ) );
DFF_X1 \myifu/myicache/_2970_ ( .D(\myifu/myicache/_1801_ ), .CK(clock ), .Q(\myifu/myicache/data[3][4] ), .QN(\myifu/myicache/_1402_ ) );
DFF_X1 \myifu/myicache/_2971_ ( .D(\myifu/myicache/_1802_ ), .CK(clock ), .Q(\myifu/myicache/data[3][5] ), .QN(\myifu/myicache/_1401_ ) );
DFF_X1 \myifu/myicache/_2972_ ( .D(\myifu/myicache/_1803_ ), .CK(clock ), .Q(\myifu/myicache/data[3][6] ), .QN(\myifu/myicache/_1400_ ) );
DFF_X1 \myifu/myicache/_2973_ ( .D(\myifu/myicache/_1804_ ), .CK(clock ), .Q(\myifu/myicache/data[3][7] ), .QN(\myifu/myicache/_1399_ ) );
DFF_X1 \myifu/myicache/_2974_ ( .D(\myifu/myicache/_1805_ ), .CK(clock ), .Q(\myifu/myicache/data[3][8] ), .QN(\myifu/myicache/_1398_ ) );
DFF_X1 \myifu/myicache/_2975_ ( .D(\myifu/myicache/_1806_ ), .CK(clock ), .Q(\myifu/myicache/data[3][9] ), .QN(\myifu/myicache/_1397_ ) );
DFF_X1 \myifu/myicache/_2976_ ( .D(\myifu/myicache/_1807_ ), .CK(clock ), .Q(\myifu/myicache/data[3][10] ), .QN(\myifu/myicache/_1396_ ) );
DFF_X1 \myifu/myicache/_2977_ ( .D(\myifu/myicache/_1808_ ), .CK(clock ), .Q(\myifu/myicache/data[3][11] ), .QN(\myifu/myicache/_1395_ ) );
DFF_X1 \myifu/myicache/_2978_ ( .D(\myifu/myicache/_1809_ ), .CK(clock ), .Q(\myifu/myicache/data[3][12] ), .QN(\myifu/myicache/_1394_ ) );
DFF_X1 \myifu/myicache/_2979_ ( .D(\myifu/myicache/_1810_ ), .CK(clock ), .Q(\myifu/myicache/data[3][13] ), .QN(\myifu/myicache/_1393_ ) );
DFF_X1 \myifu/myicache/_2980_ ( .D(\myifu/myicache/_1811_ ), .CK(clock ), .Q(\myifu/myicache/data[3][14] ), .QN(\myifu/myicache/_1392_ ) );
DFF_X1 \myifu/myicache/_2981_ ( .D(\myifu/myicache/_1812_ ), .CK(clock ), .Q(\myifu/myicache/data[3][15] ), .QN(\myifu/myicache/_1391_ ) );
DFF_X1 \myifu/myicache/_2982_ ( .D(\myifu/myicache/_1813_ ), .CK(clock ), .Q(\myifu/myicache/data[3][16] ), .QN(\myifu/myicache/_1390_ ) );
DFF_X1 \myifu/myicache/_2983_ ( .D(\myifu/myicache/_1814_ ), .CK(clock ), .Q(\myifu/myicache/data[3][17] ), .QN(\myifu/myicache/_1389_ ) );
DFF_X1 \myifu/myicache/_2984_ ( .D(\myifu/myicache/_1815_ ), .CK(clock ), .Q(\myifu/myicache/data[3][18] ), .QN(\myifu/myicache/_1388_ ) );
DFF_X1 \myifu/myicache/_2985_ ( .D(\myifu/myicache/_1816_ ), .CK(clock ), .Q(\myifu/myicache/data[3][19] ), .QN(\myifu/myicache/_1387_ ) );
DFF_X1 \myifu/myicache/_2986_ ( .D(\myifu/myicache/_1817_ ), .CK(clock ), .Q(\myifu/myicache/data[3][20] ), .QN(\myifu/myicache/_1386_ ) );
DFF_X1 \myifu/myicache/_2987_ ( .D(\myifu/myicache/_1818_ ), .CK(clock ), .Q(\myifu/myicache/data[3][21] ), .QN(\myifu/myicache/_1385_ ) );
DFF_X1 \myifu/myicache/_2988_ ( .D(\myifu/myicache/_1819_ ), .CK(clock ), .Q(\myifu/myicache/data[3][22] ), .QN(\myifu/myicache/_1384_ ) );
DFF_X1 \myifu/myicache/_2989_ ( .D(\myifu/myicache/_1820_ ), .CK(clock ), .Q(\myifu/myicache/data[3][23] ), .QN(\myifu/myicache/_1383_ ) );
DFF_X1 \myifu/myicache/_2990_ ( .D(\myifu/myicache/_1821_ ), .CK(clock ), .Q(\myifu/myicache/data[3][24] ), .QN(\myifu/myicache/_1382_ ) );
DFF_X1 \myifu/myicache/_2991_ ( .D(\myifu/myicache/_1822_ ), .CK(clock ), .Q(\myifu/myicache/data[3][25] ), .QN(\myifu/myicache/_1381_ ) );
DFF_X1 \myifu/myicache/_2992_ ( .D(\myifu/myicache/_1823_ ), .CK(clock ), .Q(\myifu/myicache/data[3][26] ), .QN(\myifu/myicache/_1380_ ) );
DFF_X1 \myifu/myicache/_2993_ ( .D(\myifu/myicache/_1824_ ), .CK(clock ), .Q(\myifu/myicache/data[3][27] ), .QN(\myifu/myicache/_1379_ ) );
DFF_X1 \myifu/myicache/_2994_ ( .D(\myifu/myicache/_1825_ ), .CK(clock ), .Q(\myifu/myicache/data[3][28] ), .QN(\myifu/myicache/_1378_ ) );
DFF_X1 \myifu/myicache/_2995_ ( .D(\myifu/myicache/_1826_ ), .CK(clock ), .Q(\myifu/myicache/data[3][29] ), .QN(\myifu/myicache/_1377_ ) );
DFF_X1 \myifu/myicache/_2996_ ( .D(\myifu/myicache/_1827_ ), .CK(clock ), .Q(\myifu/myicache/data[3][30] ), .QN(\myifu/myicache/_1376_ ) );
DFF_X1 \myifu/myicache/_2997_ ( .D(\myifu/myicache/_1828_ ), .CK(clock ), .Q(\myifu/myicache/data[3][31] ), .QN(\myifu/myicache/_1375_ ) );
DFF_X1 \myifu/myicache/_2998_ ( .D(\myifu/myicache/_1829_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][0] ), .QN(\myifu/myicache/_1374_ ) );
DFF_X1 \myifu/myicache/_2999_ ( .D(\myifu/myicache/_1830_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][1] ), .QN(\myifu/myicache/_1373_ ) );
DFF_X1 \myifu/myicache/_3000_ ( .D(\myifu/myicache/_1831_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][2] ), .QN(\myifu/myicache/_1372_ ) );
DFF_X1 \myifu/myicache/_3001_ ( .D(\myifu/myicache/_1832_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][3] ), .QN(\myifu/myicache/_1371_ ) );
DFF_X1 \myifu/myicache/_3002_ ( .D(\myifu/myicache/_1833_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][4] ), .QN(\myifu/myicache/_1370_ ) );
DFF_X1 \myifu/myicache/_3003_ ( .D(\myifu/myicache/_1834_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][5] ), .QN(\myifu/myicache/_1369_ ) );
DFF_X1 \myifu/myicache/_3004_ ( .D(\myifu/myicache/_1835_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][6] ), .QN(\myifu/myicache/_1368_ ) );
DFF_X1 \myifu/myicache/_3005_ ( .D(\myifu/myicache/_1836_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][7] ), .QN(\myifu/myicache/_1367_ ) );
DFF_X1 \myifu/myicache/_3006_ ( .D(\myifu/myicache/_1837_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][8] ), .QN(\myifu/myicache/_1366_ ) );
DFF_X1 \myifu/myicache/_3007_ ( .D(\myifu/myicache/_1838_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][9] ), .QN(\myifu/myicache/_1365_ ) );
DFF_X1 \myifu/myicache/_3008_ ( .D(\myifu/myicache/_1839_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][10] ), .QN(\myifu/myicache/_1364_ ) );
DFF_X1 \myifu/myicache/_3009_ ( .D(\myifu/myicache/_1840_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][11] ), .QN(\myifu/myicache/_1363_ ) );
DFF_X1 \myifu/myicache/_3010_ ( .D(\myifu/myicache/_1841_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][12] ), .QN(\myifu/myicache/_1362_ ) );
DFF_X1 \myifu/myicache/_3011_ ( .D(\myifu/myicache/_1842_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][13] ), .QN(\myifu/myicache/_1361_ ) );
DFF_X1 \myifu/myicache/_3012_ ( .D(\myifu/myicache/_1843_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][14] ), .QN(\myifu/myicache/_1360_ ) );
DFF_X1 \myifu/myicache/_3013_ ( .D(\myifu/myicache/_1844_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][15] ), .QN(\myifu/myicache/_1359_ ) );
DFF_X1 \myifu/myicache/_3014_ ( .D(\myifu/myicache/_1845_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][16] ), .QN(\myifu/myicache/_1358_ ) );
DFF_X1 \myifu/myicache/_3015_ ( .D(\myifu/myicache/_1846_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][17] ), .QN(\myifu/myicache/_1357_ ) );
DFF_X1 \myifu/myicache/_3016_ ( .D(\myifu/myicache/_1847_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][18] ), .QN(\myifu/myicache/_1356_ ) );
DFF_X1 \myifu/myicache/_3017_ ( .D(\myifu/myicache/_1848_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][19] ), .QN(\myifu/myicache/_1355_ ) );
DFF_X1 \myifu/myicache/_3018_ ( .D(\myifu/myicache/_1849_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][20] ), .QN(\myifu/myicache/_1354_ ) );
DFF_X1 \myifu/myicache/_3019_ ( .D(\myifu/myicache/_1850_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][21] ), .QN(\myifu/myicache/_1353_ ) );
DFF_X1 \myifu/myicache/_3020_ ( .D(\myifu/myicache/_1851_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][22] ), .QN(\myifu/myicache/_1352_ ) );
DFF_X1 \myifu/myicache/_3021_ ( .D(\myifu/myicache/_1852_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][23] ), .QN(\myifu/myicache/_1351_ ) );
DFF_X1 \myifu/myicache/_3022_ ( .D(\myifu/myicache/_1853_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][24] ), .QN(\myifu/myicache/_1350_ ) );
DFF_X1 \myifu/myicache/_3023_ ( .D(\myifu/myicache/_1854_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][25] ), .QN(\myifu/myicache/_1349_ ) );
DFF_X1 \myifu/myicache/_3024_ ( .D(\myifu/myicache/_1855_ ), .CK(clock ), .Q(\myifu/myicache/tag[2][26] ), .QN(\myifu/myicache/_1348_ ) );
DFF_X1 \myifu/myicache/_3025_ ( .D(\myifu/myicache/_1856_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][0] ), .QN(\myifu/myicache/_1347_ ) );
DFF_X1 \myifu/myicache/_3026_ ( .D(\myifu/myicache/_1857_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][1] ), .QN(\myifu/myicache/_1346_ ) );
DFF_X1 \myifu/myicache/_3027_ ( .D(\myifu/myicache/_1858_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][2] ), .QN(\myifu/myicache/_1345_ ) );
DFF_X1 \myifu/myicache/_3028_ ( .D(\myifu/myicache/_1859_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][3] ), .QN(\myifu/myicache/_1344_ ) );
DFF_X1 \myifu/myicache/_3029_ ( .D(\myifu/myicache/_1860_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][4] ), .QN(\myifu/myicache/_1343_ ) );
DFF_X1 \myifu/myicache/_3030_ ( .D(\myifu/myicache/_1861_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][5] ), .QN(\myifu/myicache/_1342_ ) );
DFF_X1 \myifu/myicache/_3031_ ( .D(\myifu/myicache/_1862_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][6] ), .QN(\myifu/myicache/_1341_ ) );
DFF_X1 \myifu/myicache/_3032_ ( .D(\myifu/myicache/_1863_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][7] ), .QN(\myifu/myicache/_1340_ ) );
DFF_X1 \myifu/myicache/_3033_ ( .D(\myifu/myicache/_1864_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][8] ), .QN(\myifu/myicache/_1339_ ) );
DFF_X1 \myifu/myicache/_3034_ ( .D(\myifu/myicache/_1865_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][9] ), .QN(\myifu/myicache/_1338_ ) );
DFF_X1 \myifu/myicache/_3035_ ( .D(\myifu/myicache/_1866_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][10] ), .QN(\myifu/myicache/_1337_ ) );
DFF_X1 \myifu/myicache/_3036_ ( .D(\myifu/myicache/_1867_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][11] ), .QN(\myifu/myicache/_1336_ ) );
DFF_X1 \myifu/myicache/_3037_ ( .D(\myifu/myicache/_1868_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][12] ), .QN(\myifu/myicache/_1335_ ) );
DFF_X1 \myifu/myicache/_3038_ ( .D(\myifu/myicache/_1869_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][13] ), .QN(\myifu/myicache/_1334_ ) );
DFF_X1 \myifu/myicache/_3039_ ( .D(\myifu/myicache/_1870_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][14] ), .QN(\myifu/myicache/_1333_ ) );
DFF_X1 \myifu/myicache/_3040_ ( .D(\myifu/myicache/_1871_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][15] ), .QN(\myifu/myicache/_1332_ ) );
DFF_X1 \myifu/myicache/_3041_ ( .D(\myifu/myicache/_1872_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][16] ), .QN(\myifu/myicache/_1331_ ) );
DFF_X1 \myifu/myicache/_3042_ ( .D(\myifu/myicache/_1873_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][17] ), .QN(\myifu/myicache/_1330_ ) );
DFF_X1 \myifu/myicache/_3043_ ( .D(\myifu/myicache/_1874_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][18] ), .QN(\myifu/myicache/_1329_ ) );
DFF_X1 \myifu/myicache/_3044_ ( .D(\myifu/myicache/_1875_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][19] ), .QN(\myifu/myicache/_1328_ ) );
DFF_X1 \myifu/myicache/_3045_ ( .D(\myifu/myicache/_1876_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][20] ), .QN(\myifu/myicache/_1327_ ) );
DFF_X1 \myifu/myicache/_3046_ ( .D(\myifu/myicache/_1877_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][21] ), .QN(\myifu/myicache/_1326_ ) );
DFF_X1 \myifu/myicache/_3047_ ( .D(\myifu/myicache/_1878_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][22] ), .QN(\myifu/myicache/_1325_ ) );
DFF_X1 \myifu/myicache/_3048_ ( .D(\myifu/myicache/_1879_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][23] ), .QN(\myifu/myicache/_1324_ ) );
DFF_X1 \myifu/myicache/_3049_ ( .D(\myifu/myicache/_1880_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][24] ), .QN(\myifu/myicache/_1323_ ) );
DFF_X1 \myifu/myicache/_3050_ ( .D(\myifu/myicache/_1881_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][25] ), .QN(\myifu/myicache/_1322_ ) );
DFF_X1 \myifu/myicache/_3051_ ( .D(\myifu/myicache/_1882_ ), .CK(clock ), .Q(\myifu/myicache/tag[1][26] ), .QN(\myifu/myicache/_1321_ ) );
DFF_X1 \myifu/myicache/_3052_ ( .D(\myifu/myicache/_1883_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][0] ), .QN(\myifu/myicache/_1320_ ) );
DFF_X1 \myifu/myicache/_3053_ ( .D(\myifu/myicache/_1884_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][1] ), .QN(\myifu/myicache/_1319_ ) );
DFF_X1 \myifu/myicache/_3054_ ( .D(\myifu/myicache/_1885_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][2] ), .QN(\myifu/myicache/_1318_ ) );
DFF_X1 \myifu/myicache/_3055_ ( .D(\myifu/myicache/_1886_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][3] ), .QN(\myifu/myicache/_1317_ ) );
DFF_X1 \myifu/myicache/_3056_ ( .D(\myifu/myicache/_1887_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][4] ), .QN(\myifu/myicache/_1316_ ) );
DFF_X1 \myifu/myicache/_3057_ ( .D(\myifu/myicache/_1888_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][5] ), .QN(\myifu/myicache/_1315_ ) );
DFF_X1 \myifu/myicache/_3058_ ( .D(\myifu/myicache/_1889_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][6] ), .QN(\myifu/myicache/_1314_ ) );
DFF_X1 \myifu/myicache/_3059_ ( .D(\myifu/myicache/_1890_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][7] ), .QN(\myifu/myicache/_1313_ ) );
DFF_X1 \myifu/myicache/_3060_ ( .D(\myifu/myicache/_1891_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][8] ), .QN(\myifu/myicache/_1312_ ) );
DFF_X1 \myifu/myicache/_3061_ ( .D(\myifu/myicache/_1892_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][9] ), .QN(\myifu/myicache/_1311_ ) );
DFF_X1 \myifu/myicache/_3062_ ( .D(\myifu/myicache/_1893_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][10] ), .QN(\myifu/myicache/_1310_ ) );
DFF_X1 \myifu/myicache/_3063_ ( .D(\myifu/myicache/_1894_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][11] ), .QN(\myifu/myicache/_1309_ ) );
DFF_X1 \myifu/myicache/_3064_ ( .D(\myifu/myicache/_1895_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][12] ), .QN(\myifu/myicache/_1308_ ) );
DFF_X1 \myifu/myicache/_3065_ ( .D(\myifu/myicache/_1896_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][13] ), .QN(\myifu/myicache/_1307_ ) );
DFF_X1 \myifu/myicache/_3066_ ( .D(\myifu/myicache/_1897_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][14] ), .QN(\myifu/myicache/_1306_ ) );
DFF_X1 \myifu/myicache/_3067_ ( .D(\myifu/myicache/_1898_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][15] ), .QN(\myifu/myicache/_1305_ ) );
DFF_X1 \myifu/myicache/_3068_ ( .D(\myifu/myicache/_1899_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][16] ), .QN(\myifu/myicache/_1304_ ) );
DFF_X1 \myifu/myicache/_3069_ ( .D(\myifu/myicache/_1900_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][17] ), .QN(\myifu/myicache/_1303_ ) );
DFF_X1 \myifu/myicache/_3070_ ( .D(\myifu/myicache/_1901_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][18] ), .QN(\myifu/myicache/_1302_ ) );
DFF_X1 \myifu/myicache/_3071_ ( .D(\myifu/myicache/_1902_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][19] ), .QN(\myifu/myicache/_1301_ ) );
DFF_X1 \myifu/myicache/_3072_ ( .D(\myifu/myicache/_1903_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][20] ), .QN(\myifu/myicache/_1300_ ) );
DFF_X1 \myifu/myicache/_3073_ ( .D(\myifu/myicache/_1904_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][21] ), .QN(\myifu/myicache/_1299_ ) );
DFF_X1 \myifu/myicache/_3074_ ( .D(\myifu/myicache/_1905_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][22] ), .QN(\myifu/myicache/_1298_ ) );
DFF_X1 \myifu/myicache/_3075_ ( .D(\myifu/myicache/_1906_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][23] ), .QN(\myifu/myicache/_1297_ ) );
DFF_X1 \myifu/myicache/_3076_ ( .D(\myifu/myicache/_1907_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][24] ), .QN(\myifu/myicache/_1296_ ) );
DFF_X1 \myifu/myicache/_3077_ ( .D(\myifu/myicache/_1908_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][25] ), .QN(\myifu/myicache/_1295_ ) );
DFF_X1 \myifu/myicache/_3078_ ( .D(\myifu/myicache/_1909_ ), .CK(clock ), .Q(\myifu/myicache/tag[0][26] ), .QN(\myifu/myicache/_1294_ ) );
DFF_X1 \myifu/myicache/_3079_ ( .D(\myifu/myicache/_1910_ ), .CK(clock ), .Q(\myifu/myicache/data[7][0] ), .QN(\myifu/myicache/_1293_ ) );
DFF_X1 \myifu/myicache/_3080_ ( .D(\myifu/myicache/_1911_ ), .CK(clock ), .Q(\myifu/myicache/data[7][1] ), .QN(\myifu/myicache/_1292_ ) );
DFF_X1 \myifu/myicache/_3081_ ( .D(\myifu/myicache/_1912_ ), .CK(clock ), .Q(\myifu/myicache/data[7][2] ), .QN(\myifu/myicache/_1291_ ) );
DFF_X1 \myifu/myicache/_3082_ ( .D(\myifu/myicache/_1913_ ), .CK(clock ), .Q(\myifu/myicache/data[7][3] ), .QN(\myifu/myicache/_1290_ ) );
DFF_X1 \myifu/myicache/_3083_ ( .D(\myifu/myicache/_1914_ ), .CK(clock ), .Q(\myifu/myicache/data[7][4] ), .QN(\myifu/myicache/_1289_ ) );
DFF_X1 \myifu/myicache/_3084_ ( .D(\myifu/myicache/_1915_ ), .CK(clock ), .Q(\myifu/myicache/data[7][5] ), .QN(\myifu/myicache/_1288_ ) );
DFF_X1 \myifu/myicache/_3085_ ( .D(\myifu/myicache/_1916_ ), .CK(clock ), .Q(\myifu/myicache/data[7][6] ), .QN(\myifu/myicache/_1287_ ) );
DFF_X1 \myifu/myicache/_3086_ ( .D(\myifu/myicache/_1917_ ), .CK(clock ), .Q(\myifu/myicache/data[7][7] ), .QN(\myifu/myicache/_1286_ ) );
DFF_X1 \myifu/myicache/_3087_ ( .D(\myifu/myicache/_1918_ ), .CK(clock ), .Q(\myifu/myicache/data[7][8] ), .QN(\myifu/myicache/_1285_ ) );
DFF_X1 \myifu/myicache/_3088_ ( .D(\myifu/myicache/_1919_ ), .CK(clock ), .Q(\myifu/myicache/data[7][9] ), .QN(\myifu/myicache/_1284_ ) );
DFF_X1 \myifu/myicache/_3089_ ( .D(\myifu/myicache/_1920_ ), .CK(clock ), .Q(\myifu/myicache/data[7][10] ), .QN(\myifu/myicache/_1283_ ) );
DFF_X1 \myifu/myicache/_3090_ ( .D(\myifu/myicache/_1921_ ), .CK(clock ), .Q(\myifu/myicache/data[7][11] ), .QN(\myifu/myicache/_1282_ ) );
DFF_X1 \myifu/myicache/_3091_ ( .D(\myifu/myicache/_1922_ ), .CK(clock ), .Q(\myifu/myicache/data[7][12] ), .QN(\myifu/myicache/_1281_ ) );
DFF_X1 \myifu/myicache/_3092_ ( .D(\myifu/myicache/_1923_ ), .CK(clock ), .Q(\myifu/myicache/data[7][13] ), .QN(\myifu/myicache/_1280_ ) );
DFF_X1 \myifu/myicache/_3093_ ( .D(\myifu/myicache/_1924_ ), .CK(clock ), .Q(\myifu/myicache/data[7][14] ), .QN(\myifu/myicache/_1279_ ) );
DFF_X1 \myifu/myicache/_3094_ ( .D(\myifu/myicache/_1925_ ), .CK(clock ), .Q(\myifu/myicache/data[7][15] ), .QN(\myifu/myicache/_1278_ ) );
DFF_X1 \myifu/myicache/_3095_ ( .D(\myifu/myicache/_1926_ ), .CK(clock ), .Q(\myifu/myicache/data[7][16] ), .QN(\myifu/myicache/_1277_ ) );
DFF_X1 \myifu/myicache/_3096_ ( .D(\myifu/myicache/_1927_ ), .CK(clock ), .Q(\myifu/myicache/data[7][17] ), .QN(\myifu/myicache/_1276_ ) );
DFF_X1 \myifu/myicache/_3097_ ( .D(\myifu/myicache/_1928_ ), .CK(clock ), .Q(\myifu/myicache/data[7][18] ), .QN(\myifu/myicache/_1275_ ) );
DFF_X1 \myifu/myicache/_3098_ ( .D(\myifu/myicache/_1929_ ), .CK(clock ), .Q(\myifu/myicache/data[7][19] ), .QN(\myifu/myicache/_1274_ ) );
DFF_X1 \myifu/myicache/_3099_ ( .D(\myifu/myicache/_1930_ ), .CK(clock ), .Q(\myifu/myicache/data[7][20] ), .QN(\myifu/myicache/_1273_ ) );
DFF_X1 \myifu/myicache/_3100_ ( .D(\myifu/myicache/_1931_ ), .CK(clock ), .Q(\myifu/myicache/data[7][21] ), .QN(\myifu/myicache/_1272_ ) );
DFF_X1 \myifu/myicache/_3101_ ( .D(\myifu/myicache/_1932_ ), .CK(clock ), .Q(\myifu/myicache/data[7][22] ), .QN(\myifu/myicache/_1271_ ) );
DFF_X1 \myifu/myicache/_3102_ ( .D(\myifu/myicache/_1933_ ), .CK(clock ), .Q(\myifu/myicache/data[7][23] ), .QN(\myifu/myicache/_1270_ ) );
DFF_X1 \myifu/myicache/_3103_ ( .D(\myifu/myicache/_1934_ ), .CK(clock ), .Q(\myifu/myicache/data[7][24] ), .QN(\myifu/myicache/_1269_ ) );
DFF_X1 \myifu/myicache/_3104_ ( .D(\myifu/myicache/_1935_ ), .CK(clock ), .Q(\myifu/myicache/data[7][25] ), .QN(\myifu/myicache/_1268_ ) );
DFF_X1 \myifu/myicache/_3105_ ( .D(\myifu/myicache/_1936_ ), .CK(clock ), .Q(\myifu/myicache/data[7][26] ), .QN(\myifu/myicache/_1267_ ) );
DFF_X1 \myifu/myicache/_3106_ ( .D(\myifu/myicache/_1937_ ), .CK(clock ), .Q(\myifu/myicache/data[7][27] ), .QN(\myifu/myicache/_1266_ ) );
DFF_X1 \myifu/myicache/_3107_ ( .D(\myifu/myicache/_1938_ ), .CK(clock ), .Q(\myifu/myicache/data[7][28] ), .QN(\myifu/myicache/_1265_ ) );
DFF_X1 \myifu/myicache/_3108_ ( .D(\myifu/myicache/_1939_ ), .CK(clock ), .Q(\myifu/myicache/data[7][29] ), .QN(\myifu/myicache/_1264_ ) );
DFF_X1 \myifu/myicache/_3109_ ( .D(\myifu/myicache/_1940_ ), .CK(clock ), .Q(\myifu/myicache/data[7][30] ), .QN(\myifu/myicache/_1263_ ) );
DFF_X1 \myifu/myicache/_3110_ ( .D(\myifu/myicache/_1941_ ), .CK(clock ), .Q(\myifu/myicache/data[7][31] ), .QN(\myifu/myicache/_1262_ ) );
DFF_X1 \myifu/myicache/_3111_ ( .D(\myifu/myicache/_1942_ ), .CK(clock ), .Q(\myifu/myicache/valid [1] ), .QN(\myifu/myicache/_1261_ ) );
DFF_X1 \myifu/myicache/_3112_ ( .D(\myifu/myicache/_1943_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][0] ), .QN(\myifu/myicache/_1260_ ) );
DFF_X1 \myifu/myicache/_3113_ ( .D(\myifu/myicache/_1944_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][1] ), .QN(\myifu/myicache/_1259_ ) );
DFF_X1 \myifu/myicache/_3114_ ( .D(\myifu/myicache/_1945_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][2] ), .QN(\myifu/myicache/_1258_ ) );
DFF_X1 \myifu/myicache/_3115_ ( .D(\myifu/myicache/_1946_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][3] ), .QN(\myifu/myicache/_1257_ ) );
DFF_X1 \myifu/myicache/_3116_ ( .D(\myifu/myicache/_1947_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][4] ), .QN(\myifu/myicache/_1256_ ) );
DFF_X1 \myifu/myicache/_3117_ ( .D(\myifu/myicache/_1948_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][5] ), .QN(\myifu/myicache/_1255_ ) );
DFF_X1 \myifu/myicache/_3118_ ( .D(\myifu/myicache/_1949_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][6] ), .QN(\myifu/myicache/_1254_ ) );
DFF_X1 \myifu/myicache/_3119_ ( .D(\myifu/myicache/_1950_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][7] ), .QN(\myifu/myicache/_1253_ ) );
DFF_X1 \myifu/myicache/_3120_ ( .D(\myifu/myicache/_1951_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][8] ), .QN(\myifu/myicache/_1252_ ) );
DFF_X1 \myifu/myicache/_3121_ ( .D(\myifu/myicache/_1952_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][9] ), .QN(\myifu/myicache/_1251_ ) );
DFF_X1 \myifu/myicache/_3122_ ( .D(\myifu/myicache/_1953_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][10] ), .QN(\myifu/myicache/_1250_ ) );
DFF_X1 \myifu/myicache/_3123_ ( .D(\myifu/myicache/_1954_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][11] ), .QN(\myifu/myicache/_1249_ ) );
DFF_X1 \myifu/myicache/_3124_ ( .D(\myifu/myicache/_1955_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][12] ), .QN(\myifu/myicache/_1248_ ) );
DFF_X1 \myifu/myicache/_3125_ ( .D(\myifu/myicache/_1956_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][13] ), .QN(\myifu/myicache/_1247_ ) );
DFF_X1 \myifu/myicache/_3126_ ( .D(\myifu/myicache/_1957_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][14] ), .QN(\myifu/myicache/_1246_ ) );
DFF_X1 \myifu/myicache/_3127_ ( .D(\myifu/myicache/_1958_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][15] ), .QN(\myifu/myicache/_1245_ ) );
DFF_X1 \myifu/myicache/_3128_ ( .D(\myifu/myicache/_1959_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][16] ), .QN(\myifu/myicache/_1244_ ) );
DFF_X1 \myifu/myicache/_3129_ ( .D(\myifu/myicache/_1960_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][17] ), .QN(\myifu/myicache/_1243_ ) );
DFF_X1 \myifu/myicache/_3130_ ( .D(\myifu/myicache/_1961_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][18] ), .QN(\myifu/myicache/_1242_ ) );
DFF_X1 \myifu/myicache/_3131_ ( .D(\myifu/myicache/_1962_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][19] ), .QN(\myifu/myicache/_1241_ ) );
DFF_X1 \myifu/myicache/_3132_ ( .D(\myifu/myicache/_1963_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][20] ), .QN(\myifu/myicache/_1240_ ) );
DFF_X1 \myifu/myicache/_3133_ ( .D(\myifu/myicache/_1964_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][21] ), .QN(\myifu/myicache/_1239_ ) );
DFF_X1 \myifu/myicache/_3134_ ( .D(\myifu/myicache/_1965_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][22] ), .QN(\myifu/myicache/_1238_ ) );
DFF_X1 \myifu/myicache/_3135_ ( .D(\myifu/myicache/_1966_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][23] ), .QN(\myifu/myicache/_1237_ ) );
DFF_X1 \myifu/myicache/_3136_ ( .D(\myifu/myicache/_1967_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][24] ), .QN(\myifu/myicache/_1236_ ) );
DFF_X1 \myifu/myicache/_3137_ ( .D(\myifu/myicache/_1968_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][25] ), .QN(\myifu/myicache/_1235_ ) );
DFF_X1 \myifu/myicache/_3138_ ( .D(\myifu/myicache/_1969_ ), .CK(clock ), .Q(\myifu/myicache/tag[3][26] ), .QN(\myifu/myicache/_1234_ ) );
BUF_X1 \myifu/myicache/_3139_ ( .A(\araddr_IFU [3] ), .Z(\myifu/myicache/_0688_ ) );
BUF_X1 \myifu/myicache/_3140_ ( .A(\araddr_IFU [4] ), .Z(\myifu/myicache/_0689_ ) );
BUF_X1 \myifu/myicache/_3141_ ( .A(\myifu/_0004_ ), .Z(\myifu/myicache/_1064_ ) );
BUF_X1 \myifu/myicache/_3142_ ( .A(\myifu/valid_in ), .Z(\myifu/myicache/_1233_ ) );
BUF_X1 \myifu/myicache/_3143_ ( .A(\myifu/offset [2] ), .Z(\myifu/myicache/_1063_ ) );
BUF_X1 \myifu/myicache/_3144_ ( .A(\myifu/valid_in ), .Z(\myifu/myicache/_1231_ ) );
BUF_X1 \myifu/myicache/_3145_ ( .A(\myifu/myicache/tag[0][0] ), .Z(\myifu/myicache/_1065_ ) );
BUF_X1 \myifu/myicache/_3146_ ( .A(\myifu/myicache/tag[1][0] ), .Z(\myifu/myicache/_1092_ ) );
BUF_X1 \myifu/myicache/_3147_ ( .A(\myifu/myicache/tag[2][0] ), .Z(\myifu/myicache/_1119_ ) );
BUF_X1 \myifu/myicache/_3148_ ( .A(\myifu/myicache/tag[3][0] ), .Z(\myifu/myicache/_1146_ ) );
BUF_X1 \myifu/myicache/_3149_ ( .A(\myifu/myicache/_1200_ ), .Z(\myifu/tag_out [0] ) );
BUF_X1 \myifu/myicache/_3150_ ( .A(\myifu/myicache/tag[0][1] ), .Z(\myifu/myicache/_1076_ ) );
BUF_X1 \myifu/myicache/_3151_ ( .A(\myifu/myicache/tag[1][1] ), .Z(\myifu/myicache/_1103_ ) );
BUF_X1 \myifu/myicache/_3152_ ( .A(\myifu/myicache/tag[2][1] ), .Z(\myifu/myicache/_1130_ ) );
BUF_X1 \myifu/myicache/_3153_ ( .A(\myifu/myicache/tag[3][1] ), .Z(\myifu/myicache/_1157_ ) );
BUF_X1 \myifu/myicache/_3154_ ( .A(\myifu/myicache/_1211_ ), .Z(\myifu/tag_out [1] ) );
BUF_X1 \myifu/myicache/_3155_ ( .A(\myifu/myicache/tag[0][2] ), .Z(\myifu/myicache/_1084_ ) );
BUF_X1 \myifu/myicache/_3156_ ( .A(\myifu/myicache/tag[1][2] ), .Z(\myifu/myicache/_1111_ ) );
BUF_X1 \myifu/myicache/_3157_ ( .A(\myifu/myicache/tag[2][2] ), .Z(\myifu/myicache/_1138_ ) );
BUF_X1 \myifu/myicache/_3158_ ( .A(\myifu/myicache/tag[3][2] ), .Z(\myifu/myicache/_1165_ ) );
BUF_X1 \myifu/myicache/_3159_ ( .A(\myifu/myicache/_1219_ ), .Z(\myifu/tag_out [2] ) );
BUF_X1 \myifu/myicache/_3160_ ( .A(\myifu/myicache/tag[0][3] ), .Z(\myifu/myicache/_1085_ ) );
BUF_X1 \myifu/myicache/_3161_ ( .A(\myifu/myicache/tag[1][3] ), .Z(\myifu/myicache/_1112_ ) );
BUF_X1 \myifu/myicache/_3162_ ( .A(\myifu/myicache/tag[2][3] ), .Z(\myifu/myicache/_1139_ ) );
BUF_X1 \myifu/myicache/_3163_ ( .A(\myifu/myicache/tag[3][3] ), .Z(\myifu/myicache/_1166_ ) );
BUF_X1 \myifu/myicache/_3164_ ( .A(\myifu/myicache/_1220_ ), .Z(\myifu/tag_out [3] ) );
BUF_X1 \myifu/myicache/_3165_ ( .A(\myifu/myicache/tag[0][4] ), .Z(\myifu/myicache/_1086_ ) );
BUF_X1 \myifu/myicache/_3166_ ( .A(\myifu/myicache/tag[1][4] ), .Z(\myifu/myicache/_1113_ ) );
BUF_X1 \myifu/myicache/_3167_ ( .A(\myifu/myicache/tag[2][4] ), .Z(\myifu/myicache/_1140_ ) );
BUF_X1 \myifu/myicache/_3168_ ( .A(\myifu/myicache/tag[3][4] ), .Z(\myifu/myicache/_1167_ ) );
BUF_X1 \myifu/myicache/_3169_ ( .A(\myifu/myicache/_1221_ ), .Z(\myifu/tag_out [4] ) );
BUF_X1 \myifu/myicache/_3170_ ( .A(\myifu/myicache/tag[0][5] ), .Z(\myifu/myicache/_1087_ ) );
BUF_X1 \myifu/myicache/_3171_ ( .A(\myifu/myicache/tag[1][5] ), .Z(\myifu/myicache/_1114_ ) );
BUF_X1 \myifu/myicache/_3172_ ( .A(\myifu/myicache/tag[2][5] ), .Z(\myifu/myicache/_1141_ ) );
BUF_X1 \myifu/myicache/_3173_ ( .A(\myifu/myicache/tag[3][5] ), .Z(\myifu/myicache/_1168_ ) );
BUF_X1 \myifu/myicache/_3174_ ( .A(\myifu/myicache/_1222_ ), .Z(\myifu/tag_out [5] ) );
BUF_X1 \myifu/myicache/_3175_ ( .A(\myifu/myicache/tag[0][6] ), .Z(\myifu/myicache/_1088_ ) );
BUF_X1 \myifu/myicache/_3176_ ( .A(\myifu/myicache/tag[1][6] ), .Z(\myifu/myicache/_1115_ ) );
BUF_X1 \myifu/myicache/_3177_ ( .A(\myifu/myicache/tag[2][6] ), .Z(\myifu/myicache/_1142_ ) );
BUF_X1 \myifu/myicache/_3178_ ( .A(\myifu/myicache/tag[3][6] ), .Z(\myifu/myicache/_1169_ ) );
BUF_X1 \myifu/myicache/_3179_ ( .A(\myifu/myicache/_1223_ ), .Z(\myifu/tag_out [6] ) );
BUF_X1 \myifu/myicache/_3180_ ( .A(\myifu/myicache/tag[0][7] ), .Z(\myifu/myicache/_1089_ ) );
BUF_X1 \myifu/myicache/_3181_ ( .A(\myifu/myicache/tag[1][7] ), .Z(\myifu/myicache/_1116_ ) );
BUF_X1 \myifu/myicache/_3182_ ( .A(\myifu/myicache/tag[2][7] ), .Z(\myifu/myicache/_1143_ ) );
BUF_X1 \myifu/myicache/_3183_ ( .A(\myifu/myicache/tag[3][7] ), .Z(\myifu/myicache/_1170_ ) );
BUF_X1 \myifu/myicache/_3184_ ( .A(\myifu/myicache/_1224_ ), .Z(\myifu/tag_out [7] ) );
BUF_X1 \myifu/myicache/_3185_ ( .A(\myifu/myicache/tag[0][8] ), .Z(\myifu/myicache/_1090_ ) );
BUF_X1 \myifu/myicache/_3186_ ( .A(\myifu/myicache/tag[1][8] ), .Z(\myifu/myicache/_1117_ ) );
BUF_X1 \myifu/myicache/_3187_ ( .A(\myifu/myicache/tag[2][8] ), .Z(\myifu/myicache/_1144_ ) );
BUF_X1 \myifu/myicache/_3188_ ( .A(\myifu/myicache/tag[3][8] ), .Z(\myifu/myicache/_1171_ ) );
BUF_X1 \myifu/myicache/_3189_ ( .A(\myifu/myicache/_1225_ ), .Z(\myifu/tag_out [8] ) );
BUF_X1 \myifu/myicache/_3190_ ( .A(\myifu/myicache/tag[0][9] ), .Z(\myifu/myicache/_1091_ ) );
BUF_X1 \myifu/myicache/_3191_ ( .A(\myifu/myicache/tag[1][9] ), .Z(\myifu/myicache/_1118_ ) );
BUF_X1 \myifu/myicache/_3192_ ( .A(\myifu/myicache/tag[2][9] ), .Z(\myifu/myicache/_1145_ ) );
BUF_X1 \myifu/myicache/_3193_ ( .A(\myifu/myicache/tag[3][9] ), .Z(\myifu/myicache/_1172_ ) );
BUF_X1 \myifu/myicache/_3194_ ( .A(\myifu/myicache/_1226_ ), .Z(\myifu/tag_out [9] ) );
BUF_X1 \myifu/myicache/_3195_ ( .A(\myifu/myicache/tag[0][10] ), .Z(\myifu/myicache/_1066_ ) );
BUF_X1 \myifu/myicache/_3196_ ( .A(\myifu/myicache/tag[1][10] ), .Z(\myifu/myicache/_1093_ ) );
BUF_X1 \myifu/myicache/_3197_ ( .A(\myifu/myicache/tag[2][10] ), .Z(\myifu/myicache/_1120_ ) );
BUF_X1 \myifu/myicache/_3198_ ( .A(\myifu/myicache/tag[3][10] ), .Z(\myifu/myicache/_1147_ ) );
BUF_X1 \myifu/myicache/_3199_ ( .A(\myifu/myicache/_1201_ ), .Z(\myifu/tag_out [10] ) );
BUF_X1 \myifu/myicache/_3200_ ( .A(\myifu/myicache/tag[0][11] ), .Z(\myifu/myicache/_1067_ ) );
BUF_X1 \myifu/myicache/_3201_ ( .A(\myifu/myicache/tag[1][11] ), .Z(\myifu/myicache/_1094_ ) );
BUF_X1 \myifu/myicache/_3202_ ( .A(\myifu/myicache/tag[2][11] ), .Z(\myifu/myicache/_1121_ ) );
BUF_X1 \myifu/myicache/_3203_ ( .A(\myifu/myicache/tag[3][11] ), .Z(\myifu/myicache/_1148_ ) );
BUF_X1 \myifu/myicache/_3204_ ( .A(\myifu/myicache/_1202_ ), .Z(\myifu/tag_out [11] ) );
BUF_X1 \myifu/myicache/_3205_ ( .A(\myifu/myicache/tag[0][12] ), .Z(\myifu/myicache/_1068_ ) );
BUF_X1 \myifu/myicache/_3206_ ( .A(\myifu/myicache/tag[1][12] ), .Z(\myifu/myicache/_1095_ ) );
BUF_X1 \myifu/myicache/_3207_ ( .A(\myifu/myicache/tag[2][12] ), .Z(\myifu/myicache/_1122_ ) );
BUF_X1 \myifu/myicache/_3208_ ( .A(\myifu/myicache/tag[3][12] ), .Z(\myifu/myicache/_1149_ ) );
BUF_X1 \myifu/myicache/_3209_ ( .A(\myifu/myicache/_1203_ ), .Z(\myifu/tag_out [12] ) );
BUF_X1 \myifu/myicache/_3210_ ( .A(\myifu/myicache/tag[0][13] ), .Z(\myifu/myicache/_1069_ ) );
BUF_X1 \myifu/myicache/_3211_ ( .A(\myifu/myicache/tag[1][13] ), .Z(\myifu/myicache/_1096_ ) );
BUF_X1 \myifu/myicache/_3212_ ( .A(\myifu/myicache/tag[2][13] ), .Z(\myifu/myicache/_1123_ ) );
BUF_X1 \myifu/myicache/_3213_ ( .A(\myifu/myicache/tag[3][13] ), .Z(\myifu/myicache/_1150_ ) );
BUF_X1 \myifu/myicache/_3214_ ( .A(\myifu/myicache/_1204_ ), .Z(\myifu/tag_out [13] ) );
BUF_X1 \myifu/myicache/_3215_ ( .A(\myifu/myicache/tag[0][14] ), .Z(\myifu/myicache/_1070_ ) );
BUF_X1 \myifu/myicache/_3216_ ( .A(\myifu/myicache/tag[1][14] ), .Z(\myifu/myicache/_1097_ ) );
BUF_X1 \myifu/myicache/_3217_ ( .A(\myifu/myicache/tag[2][14] ), .Z(\myifu/myicache/_1124_ ) );
BUF_X1 \myifu/myicache/_3218_ ( .A(\myifu/myicache/tag[3][14] ), .Z(\myifu/myicache/_1151_ ) );
BUF_X1 \myifu/myicache/_3219_ ( .A(\myifu/myicache/_1205_ ), .Z(\myifu/tag_out [14] ) );
BUF_X1 \myifu/myicache/_3220_ ( .A(\myifu/myicache/tag[0][15] ), .Z(\myifu/myicache/_1071_ ) );
BUF_X1 \myifu/myicache/_3221_ ( .A(\myifu/myicache/tag[1][15] ), .Z(\myifu/myicache/_1098_ ) );
BUF_X1 \myifu/myicache/_3222_ ( .A(\myifu/myicache/tag[2][15] ), .Z(\myifu/myicache/_1125_ ) );
BUF_X1 \myifu/myicache/_3223_ ( .A(\myifu/myicache/tag[3][15] ), .Z(\myifu/myicache/_1152_ ) );
BUF_X1 \myifu/myicache/_3224_ ( .A(\myifu/myicache/_1206_ ), .Z(\myifu/tag_out [15] ) );
BUF_X1 \myifu/myicache/_3225_ ( .A(\myifu/myicache/tag[0][16] ), .Z(\myifu/myicache/_1072_ ) );
BUF_X1 \myifu/myicache/_3226_ ( .A(\myifu/myicache/tag[1][16] ), .Z(\myifu/myicache/_1099_ ) );
BUF_X1 \myifu/myicache/_3227_ ( .A(\myifu/myicache/tag[2][16] ), .Z(\myifu/myicache/_1126_ ) );
BUF_X1 \myifu/myicache/_3228_ ( .A(\myifu/myicache/tag[3][16] ), .Z(\myifu/myicache/_1153_ ) );
BUF_X1 \myifu/myicache/_3229_ ( .A(\myifu/myicache/_1207_ ), .Z(\myifu/tag_out [16] ) );
BUF_X1 \myifu/myicache/_3230_ ( .A(\myifu/myicache/tag[0][17] ), .Z(\myifu/myicache/_1073_ ) );
BUF_X1 \myifu/myicache/_3231_ ( .A(\myifu/myicache/tag[1][17] ), .Z(\myifu/myicache/_1100_ ) );
BUF_X1 \myifu/myicache/_3232_ ( .A(\myifu/myicache/tag[2][17] ), .Z(\myifu/myicache/_1127_ ) );
BUF_X1 \myifu/myicache/_3233_ ( .A(\myifu/myicache/tag[3][17] ), .Z(\myifu/myicache/_1154_ ) );
BUF_X1 \myifu/myicache/_3234_ ( .A(\myifu/myicache/_1208_ ), .Z(\myifu/tag_out [17] ) );
BUF_X1 \myifu/myicache/_3235_ ( .A(\myifu/myicache/tag[0][18] ), .Z(\myifu/myicache/_1074_ ) );
BUF_X1 \myifu/myicache/_3236_ ( .A(\myifu/myicache/tag[1][18] ), .Z(\myifu/myicache/_1101_ ) );
BUF_X1 \myifu/myicache/_3237_ ( .A(\myifu/myicache/tag[2][18] ), .Z(\myifu/myicache/_1128_ ) );
BUF_X1 \myifu/myicache/_3238_ ( .A(\myifu/myicache/tag[3][18] ), .Z(\myifu/myicache/_1155_ ) );
BUF_X1 \myifu/myicache/_3239_ ( .A(\myifu/myicache/_1209_ ), .Z(\myifu/tag_out [18] ) );
BUF_X1 \myifu/myicache/_3240_ ( .A(\myifu/myicache/tag[0][19] ), .Z(\myifu/myicache/_1075_ ) );
BUF_X1 \myifu/myicache/_3241_ ( .A(\myifu/myicache/tag[1][19] ), .Z(\myifu/myicache/_1102_ ) );
BUF_X1 \myifu/myicache/_3242_ ( .A(\myifu/myicache/tag[2][19] ), .Z(\myifu/myicache/_1129_ ) );
BUF_X1 \myifu/myicache/_3243_ ( .A(\myifu/myicache/tag[3][19] ), .Z(\myifu/myicache/_1156_ ) );
BUF_X1 \myifu/myicache/_3244_ ( .A(\myifu/myicache/_1210_ ), .Z(\myifu/tag_out [19] ) );
BUF_X1 \myifu/myicache/_3245_ ( .A(\myifu/myicache/tag[0][20] ), .Z(\myifu/myicache/_1077_ ) );
BUF_X1 \myifu/myicache/_3246_ ( .A(\myifu/myicache/tag[1][20] ), .Z(\myifu/myicache/_1104_ ) );
BUF_X1 \myifu/myicache/_3247_ ( .A(\myifu/myicache/tag[2][20] ), .Z(\myifu/myicache/_1131_ ) );
BUF_X1 \myifu/myicache/_3248_ ( .A(\myifu/myicache/tag[3][20] ), .Z(\myifu/myicache/_1158_ ) );
BUF_X1 \myifu/myicache/_3249_ ( .A(\myifu/myicache/_1212_ ), .Z(\myifu/tag_out [20] ) );
BUF_X1 \myifu/myicache/_3250_ ( .A(\myifu/myicache/tag[0][21] ), .Z(\myifu/myicache/_1078_ ) );
BUF_X1 \myifu/myicache/_3251_ ( .A(\myifu/myicache/tag[1][21] ), .Z(\myifu/myicache/_1105_ ) );
BUF_X1 \myifu/myicache/_3252_ ( .A(\myifu/myicache/tag[2][21] ), .Z(\myifu/myicache/_1132_ ) );
BUF_X1 \myifu/myicache/_3253_ ( .A(\myifu/myicache/tag[3][21] ), .Z(\myifu/myicache/_1159_ ) );
BUF_X1 \myifu/myicache/_3254_ ( .A(\myifu/myicache/_1213_ ), .Z(\myifu/tag_out [21] ) );
BUF_X1 \myifu/myicache/_3255_ ( .A(\myifu/myicache/tag[0][22] ), .Z(\myifu/myicache/_1079_ ) );
BUF_X1 \myifu/myicache/_3256_ ( .A(\myifu/myicache/tag[1][22] ), .Z(\myifu/myicache/_1106_ ) );
BUF_X1 \myifu/myicache/_3257_ ( .A(\myifu/myicache/tag[2][22] ), .Z(\myifu/myicache/_1133_ ) );
BUF_X1 \myifu/myicache/_3258_ ( .A(\myifu/myicache/tag[3][22] ), .Z(\myifu/myicache/_1160_ ) );
BUF_X1 \myifu/myicache/_3259_ ( .A(\myifu/myicache/_1214_ ), .Z(\myifu/tag_out [22] ) );
BUF_X1 \myifu/myicache/_3260_ ( .A(\myifu/myicache/tag[0][23] ), .Z(\myifu/myicache/_1080_ ) );
BUF_X1 \myifu/myicache/_3261_ ( .A(\myifu/myicache/tag[1][23] ), .Z(\myifu/myicache/_1107_ ) );
BUF_X1 \myifu/myicache/_3262_ ( .A(\myifu/myicache/tag[2][23] ), .Z(\myifu/myicache/_1134_ ) );
BUF_X1 \myifu/myicache/_3263_ ( .A(\myifu/myicache/tag[3][23] ), .Z(\myifu/myicache/_1161_ ) );
BUF_X1 \myifu/myicache/_3264_ ( .A(\myifu/myicache/_1215_ ), .Z(\myifu/tag_out [23] ) );
BUF_X1 \myifu/myicache/_3265_ ( .A(\myifu/myicache/tag[0][24] ), .Z(\myifu/myicache/_1081_ ) );
BUF_X1 \myifu/myicache/_3266_ ( .A(\myifu/myicache/tag[1][24] ), .Z(\myifu/myicache/_1108_ ) );
BUF_X1 \myifu/myicache/_3267_ ( .A(\myifu/myicache/tag[2][24] ), .Z(\myifu/myicache/_1135_ ) );
BUF_X1 \myifu/myicache/_3268_ ( .A(\myifu/myicache/tag[3][24] ), .Z(\myifu/myicache/_1162_ ) );
BUF_X1 \myifu/myicache/_3269_ ( .A(\myifu/myicache/_1216_ ), .Z(\myifu/tag_out [24] ) );
BUF_X1 \myifu/myicache/_3270_ ( .A(\myifu/myicache/tag[0][25] ), .Z(\myifu/myicache/_1082_ ) );
BUF_X1 \myifu/myicache/_3271_ ( .A(\myifu/myicache/tag[1][25] ), .Z(\myifu/myicache/_1109_ ) );
BUF_X1 \myifu/myicache/_3272_ ( .A(\myifu/myicache/tag[2][25] ), .Z(\myifu/myicache/_1136_ ) );
BUF_X1 \myifu/myicache/_3273_ ( .A(\myifu/myicache/tag[3][25] ), .Z(\myifu/myicache/_1163_ ) );
BUF_X1 \myifu/myicache/_3274_ ( .A(\myifu/myicache/_1217_ ), .Z(\myifu/tag_out [25] ) );
BUF_X1 \myifu/myicache/_3275_ ( .A(\myifu/myicache/tag[0][26] ), .Z(\myifu/myicache/_1083_ ) );
BUF_X1 \myifu/myicache/_3276_ ( .A(\myifu/myicache/tag[1][26] ), .Z(\myifu/myicache/_1110_ ) );
BUF_X1 \myifu/myicache/_3277_ ( .A(\myifu/myicache/tag[2][26] ), .Z(\myifu/myicache/_1137_ ) );
BUF_X1 \myifu/myicache/_3278_ ( .A(\myifu/myicache/tag[3][26] ), .Z(\myifu/myicache/_1164_ ) );
BUF_X1 \myifu/myicache/_3279_ ( .A(\myifu/myicache/_1218_ ), .Z(\myifu/tag_out [26] ) );
BUF_X1 \myifu/myicache/_3280_ ( .A(\myifu/myicache/valid [0] ), .Z(\myifu/myicache/_1227_ ) );
BUF_X1 \myifu/myicache/_3281_ ( .A(\myifu/myicache/valid [1] ), .Z(\myifu/myicache/_1228_ ) );
BUF_X1 \myifu/myicache/_3282_ ( .A(\myifu/myicache/valid [2] ), .Z(\myifu/myicache/_1229_ ) );
BUF_X1 \myifu/myicache/_3283_ ( .A(\myifu/myicache/valid [3] ), .Z(\myifu/myicache/_1230_ ) );
BUF_X1 \myifu/myicache/_3284_ ( .A(\myifu/myicache/_1232_ ), .Z(\myifu/valid_out ) );
BUF_X1 \myifu/myicache/_3285_ ( .A(\myifu/myicache/data[0][0] ), .Z(\myifu/myicache/_0368_ ) );
BUF_X1 \myifu/myicache/_3286_ ( .A(\myifu/myicache/data[1][0] ), .Z(\myifu/myicache/_0400_ ) );
BUF_X1 \myifu/myicache/_3287_ ( .A(\myifu/myicache/data[2][0] ), .Z(\myifu/myicache/_0432_ ) );
BUF_X1 \myifu/myicache/_3288_ ( .A(\myifu/myicache/data[3][0] ), .Z(\myifu/myicache/_0464_ ) );
BUF_X1 \myifu/myicache/_3289_ ( .A(\myifu/myicache/data[4][0] ), .Z(\myifu/myicache/_0496_ ) );
BUF_X1 \myifu/myicache/_3290_ ( .A(\myifu/myicache/data[5][0] ), .Z(\myifu/myicache/_0528_ ) );
BUF_X1 \myifu/myicache/_3291_ ( .A(\myifu/myicache/data[6][0] ), .Z(\myifu/myicache/_0560_ ) );
BUF_X1 \myifu/myicache/_3292_ ( .A(\myifu/myicache/data[7][0] ), .Z(\myifu/myicache/_0592_ ) );
BUF_X1 \myifu/myicache/_3293_ ( .A(\myifu/myicache/_0656_ ), .Z(\myifu/data_out [0] ) );
BUF_X1 \myifu/myicache/_3294_ ( .A(\myifu/myicache/data[0][1] ), .Z(\myifu/myicache/_0379_ ) );
BUF_X1 \myifu/myicache/_3295_ ( .A(\myifu/myicache/data[1][1] ), .Z(\myifu/myicache/_0411_ ) );
BUF_X1 \myifu/myicache/_3296_ ( .A(\myifu/myicache/data[2][1] ), .Z(\myifu/myicache/_0443_ ) );
BUF_X1 \myifu/myicache/_3297_ ( .A(\myifu/myicache/data[3][1] ), .Z(\myifu/myicache/_0475_ ) );
BUF_X1 \myifu/myicache/_3298_ ( .A(\myifu/myicache/data[4][1] ), .Z(\myifu/myicache/_0507_ ) );
BUF_X1 \myifu/myicache/_3299_ ( .A(\myifu/myicache/data[5][1] ), .Z(\myifu/myicache/_0539_ ) );
BUF_X1 \myifu/myicache/_3300_ ( .A(\myifu/myicache/data[6][1] ), .Z(\myifu/myicache/_0571_ ) );
BUF_X1 \myifu/myicache/_3301_ ( .A(\myifu/myicache/data[7][1] ), .Z(\myifu/myicache/_0603_ ) );
BUF_X1 \myifu/myicache/_3302_ ( .A(\myifu/myicache/_0667_ ), .Z(\myifu/data_out [1] ) );
BUF_X1 \myifu/myicache/_3303_ ( .A(\myifu/myicache/data[0][2] ), .Z(\myifu/myicache/_0390_ ) );
BUF_X1 \myifu/myicache/_3304_ ( .A(\myifu/myicache/data[1][2] ), .Z(\myifu/myicache/_0422_ ) );
BUF_X1 \myifu/myicache/_3305_ ( .A(\myifu/myicache/data[2][2] ), .Z(\myifu/myicache/_0454_ ) );
BUF_X1 \myifu/myicache/_3306_ ( .A(\myifu/myicache/data[3][2] ), .Z(\myifu/myicache/_0486_ ) );
BUF_X1 \myifu/myicache/_3307_ ( .A(\myifu/myicache/data[4][2] ), .Z(\myifu/myicache/_0518_ ) );
BUF_X1 \myifu/myicache/_3308_ ( .A(\myifu/myicache/data[5][2] ), .Z(\myifu/myicache/_0550_ ) );
BUF_X1 \myifu/myicache/_3309_ ( .A(\myifu/myicache/data[6][2] ), .Z(\myifu/myicache/_0582_ ) );
BUF_X1 \myifu/myicache/_3310_ ( .A(\myifu/myicache/data[7][2] ), .Z(\myifu/myicache/_0614_ ) );
BUF_X1 \myifu/myicache/_3311_ ( .A(\myifu/myicache/_0678_ ), .Z(\myifu/data_out [2] ) );
BUF_X1 \myifu/myicache/_3312_ ( .A(\myifu/myicache/data[0][3] ), .Z(\myifu/myicache/_0393_ ) );
BUF_X1 \myifu/myicache/_3313_ ( .A(\myifu/myicache/data[1][3] ), .Z(\myifu/myicache/_0425_ ) );
BUF_X1 \myifu/myicache/_3314_ ( .A(\myifu/myicache/data[2][3] ), .Z(\myifu/myicache/_0457_ ) );
BUF_X1 \myifu/myicache/_3315_ ( .A(\myifu/myicache/data[3][3] ), .Z(\myifu/myicache/_0489_ ) );
BUF_X1 \myifu/myicache/_3316_ ( .A(\myifu/myicache/data[4][3] ), .Z(\myifu/myicache/_0521_ ) );
BUF_X1 \myifu/myicache/_3317_ ( .A(\myifu/myicache/data[5][3] ), .Z(\myifu/myicache/_0553_ ) );
BUF_X1 \myifu/myicache/_3318_ ( .A(\myifu/myicache/data[6][3] ), .Z(\myifu/myicache/_0585_ ) );
BUF_X1 \myifu/myicache/_3319_ ( .A(\myifu/myicache/data[7][3] ), .Z(\myifu/myicache/_0617_ ) );
BUF_X1 \myifu/myicache/_3320_ ( .A(\myifu/myicache/_0681_ ), .Z(\myifu/data_out [3] ) );
BUF_X1 \myifu/myicache/_3321_ ( .A(\myifu/myicache/data[0][4] ), .Z(\myifu/myicache/_0394_ ) );
BUF_X1 \myifu/myicache/_3322_ ( .A(\myifu/myicache/data[1][4] ), .Z(\myifu/myicache/_0426_ ) );
BUF_X1 \myifu/myicache/_3323_ ( .A(\myifu/myicache/data[2][4] ), .Z(\myifu/myicache/_0458_ ) );
BUF_X1 \myifu/myicache/_3324_ ( .A(\myifu/myicache/data[3][4] ), .Z(\myifu/myicache/_0490_ ) );
BUF_X1 \myifu/myicache/_3325_ ( .A(\myifu/myicache/data[4][4] ), .Z(\myifu/myicache/_0522_ ) );
BUF_X1 \myifu/myicache/_3326_ ( .A(\myifu/myicache/data[5][4] ), .Z(\myifu/myicache/_0554_ ) );
BUF_X1 \myifu/myicache/_3327_ ( .A(\myifu/myicache/data[6][4] ), .Z(\myifu/myicache/_0586_ ) );
BUF_X1 \myifu/myicache/_3328_ ( .A(\myifu/myicache/data[7][4] ), .Z(\myifu/myicache/_0618_ ) );
BUF_X1 \myifu/myicache/_3329_ ( .A(\myifu/myicache/_0682_ ), .Z(\myifu/data_out [4] ) );
BUF_X1 \myifu/myicache/_3330_ ( .A(\myifu/myicache/data[0][5] ), .Z(\myifu/myicache/_0395_ ) );
BUF_X1 \myifu/myicache/_3331_ ( .A(\myifu/myicache/data[1][5] ), .Z(\myifu/myicache/_0427_ ) );
BUF_X1 \myifu/myicache/_3332_ ( .A(\myifu/myicache/data[2][5] ), .Z(\myifu/myicache/_0459_ ) );
BUF_X1 \myifu/myicache/_3333_ ( .A(\myifu/myicache/data[3][5] ), .Z(\myifu/myicache/_0491_ ) );
BUF_X1 \myifu/myicache/_3334_ ( .A(\myifu/myicache/data[4][5] ), .Z(\myifu/myicache/_0523_ ) );
BUF_X1 \myifu/myicache/_3335_ ( .A(\myifu/myicache/data[5][5] ), .Z(\myifu/myicache/_0555_ ) );
BUF_X1 \myifu/myicache/_3336_ ( .A(\myifu/myicache/data[6][5] ), .Z(\myifu/myicache/_0587_ ) );
BUF_X1 \myifu/myicache/_3337_ ( .A(\myifu/myicache/data[7][5] ), .Z(\myifu/myicache/_0619_ ) );
BUF_X1 \myifu/myicache/_3338_ ( .A(\myifu/myicache/_0683_ ), .Z(\myifu/data_out [5] ) );
BUF_X1 \myifu/myicache/_3339_ ( .A(\myifu/myicache/data[0][6] ), .Z(\myifu/myicache/_0396_ ) );
BUF_X1 \myifu/myicache/_3340_ ( .A(\myifu/myicache/data[1][6] ), .Z(\myifu/myicache/_0428_ ) );
BUF_X1 \myifu/myicache/_3341_ ( .A(\myifu/myicache/data[2][6] ), .Z(\myifu/myicache/_0460_ ) );
BUF_X1 \myifu/myicache/_3342_ ( .A(\myifu/myicache/data[3][6] ), .Z(\myifu/myicache/_0492_ ) );
BUF_X1 \myifu/myicache/_3343_ ( .A(\myifu/myicache/data[4][6] ), .Z(\myifu/myicache/_0524_ ) );
BUF_X1 \myifu/myicache/_3344_ ( .A(\myifu/myicache/data[5][6] ), .Z(\myifu/myicache/_0556_ ) );
BUF_X1 \myifu/myicache/_3345_ ( .A(\myifu/myicache/data[6][6] ), .Z(\myifu/myicache/_0588_ ) );
BUF_X1 \myifu/myicache/_3346_ ( .A(\myifu/myicache/data[7][6] ), .Z(\myifu/myicache/_0620_ ) );
BUF_X1 \myifu/myicache/_3347_ ( .A(\myifu/myicache/_0684_ ), .Z(\myifu/data_out [6] ) );
BUF_X1 \myifu/myicache/_3348_ ( .A(\myifu/myicache/data[0][7] ), .Z(\myifu/myicache/_0397_ ) );
BUF_X1 \myifu/myicache/_3349_ ( .A(\myifu/myicache/data[1][7] ), .Z(\myifu/myicache/_0429_ ) );
BUF_X1 \myifu/myicache/_3350_ ( .A(\myifu/myicache/data[2][7] ), .Z(\myifu/myicache/_0461_ ) );
BUF_X1 \myifu/myicache/_3351_ ( .A(\myifu/myicache/data[3][7] ), .Z(\myifu/myicache/_0493_ ) );
BUF_X1 \myifu/myicache/_3352_ ( .A(\myifu/myicache/data[4][7] ), .Z(\myifu/myicache/_0525_ ) );
BUF_X1 \myifu/myicache/_3353_ ( .A(\myifu/myicache/data[5][7] ), .Z(\myifu/myicache/_0557_ ) );
BUF_X1 \myifu/myicache/_3354_ ( .A(\myifu/myicache/data[6][7] ), .Z(\myifu/myicache/_0589_ ) );
BUF_X1 \myifu/myicache/_3355_ ( .A(\myifu/myicache/data[7][7] ), .Z(\myifu/myicache/_0621_ ) );
BUF_X1 \myifu/myicache/_3356_ ( .A(\myifu/myicache/_0685_ ), .Z(\myifu/data_out [7] ) );
BUF_X1 \myifu/myicache/_3357_ ( .A(\myifu/myicache/data[0][8] ), .Z(\myifu/myicache/_0398_ ) );
BUF_X1 \myifu/myicache/_3358_ ( .A(\myifu/myicache/data[1][8] ), .Z(\myifu/myicache/_0430_ ) );
BUF_X1 \myifu/myicache/_3359_ ( .A(\myifu/myicache/data[2][8] ), .Z(\myifu/myicache/_0462_ ) );
BUF_X1 \myifu/myicache/_3360_ ( .A(\myifu/myicache/data[3][8] ), .Z(\myifu/myicache/_0494_ ) );
BUF_X1 \myifu/myicache/_3361_ ( .A(\myifu/myicache/data[4][8] ), .Z(\myifu/myicache/_0526_ ) );
BUF_X1 \myifu/myicache/_3362_ ( .A(\myifu/myicache/data[5][8] ), .Z(\myifu/myicache/_0558_ ) );
BUF_X1 \myifu/myicache/_3363_ ( .A(\myifu/myicache/data[6][8] ), .Z(\myifu/myicache/_0590_ ) );
BUF_X1 \myifu/myicache/_3364_ ( .A(\myifu/myicache/data[7][8] ), .Z(\myifu/myicache/_0622_ ) );
BUF_X1 \myifu/myicache/_3365_ ( .A(\myifu/myicache/_0686_ ), .Z(\myifu/data_out [8] ) );
BUF_X1 \myifu/myicache/_3366_ ( .A(\myifu/myicache/data[0][9] ), .Z(\myifu/myicache/_0399_ ) );
BUF_X1 \myifu/myicache/_3367_ ( .A(\myifu/myicache/data[1][9] ), .Z(\myifu/myicache/_0431_ ) );
BUF_X1 \myifu/myicache/_3368_ ( .A(\myifu/myicache/data[2][9] ), .Z(\myifu/myicache/_0463_ ) );
BUF_X1 \myifu/myicache/_3369_ ( .A(\myifu/myicache/data[3][9] ), .Z(\myifu/myicache/_0495_ ) );
BUF_X1 \myifu/myicache/_3370_ ( .A(\myifu/myicache/data[4][9] ), .Z(\myifu/myicache/_0527_ ) );
BUF_X1 \myifu/myicache/_3371_ ( .A(\myifu/myicache/data[5][9] ), .Z(\myifu/myicache/_0559_ ) );
BUF_X1 \myifu/myicache/_3372_ ( .A(\myifu/myicache/data[6][9] ), .Z(\myifu/myicache/_0591_ ) );
BUF_X1 \myifu/myicache/_3373_ ( .A(\myifu/myicache/data[7][9] ), .Z(\myifu/myicache/_0623_ ) );
BUF_X1 \myifu/myicache/_3374_ ( .A(\myifu/myicache/_0687_ ), .Z(\myifu/data_out [9] ) );
BUF_X1 \myifu/myicache/_3375_ ( .A(\myifu/myicache/data[0][10] ), .Z(\myifu/myicache/_0369_ ) );
BUF_X1 \myifu/myicache/_3376_ ( .A(\myifu/myicache/data[1][10] ), .Z(\myifu/myicache/_0401_ ) );
BUF_X1 \myifu/myicache/_3377_ ( .A(\myifu/myicache/data[2][10] ), .Z(\myifu/myicache/_0433_ ) );
BUF_X1 \myifu/myicache/_3378_ ( .A(\myifu/myicache/data[3][10] ), .Z(\myifu/myicache/_0465_ ) );
BUF_X1 \myifu/myicache/_3379_ ( .A(\myifu/myicache/data[4][10] ), .Z(\myifu/myicache/_0497_ ) );
BUF_X1 \myifu/myicache/_3380_ ( .A(\myifu/myicache/data[5][10] ), .Z(\myifu/myicache/_0529_ ) );
BUF_X1 \myifu/myicache/_3381_ ( .A(\myifu/myicache/data[6][10] ), .Z(\myifu/myicache/_0561_ ) );
BUF_X1 \myifu/myicache/_3382_ ( .A(\myifu/myicache/data[7][10] ), .Z(\myifu/myicache/_0593_ ) );
BUF_X1 \myifu/myicache/_3383_ ( .A(\myifu/myicache/_0657_ ), .Z(\myifu/data_out [10] ) );
BUF_X1 \myifu/myicache/_3384_ ( .A(\myifu/myicache/data[0][11] ), .Z(\myifu/myicache/_0370_ ) );
BUF_X1 \myifu/myicache/_3385_ ( .A(\myifu/myicache/data[1][11] ), .Z(\myifu/myicache/_0402_ ) );
BUF_X1 \myifu/myicache/_3386_ ( .A(\myifu/myicache/data[2][11] ), .Z(\myifu/myicache/_0434_ ) );
BUF_X1 \myifu/myicache/_3387_ ( .A(\myifu/myicache/data[3][11] ), .Z(\myifu/myicache/_0466_ ) );
BUF_X1 \myifu/myicache/_3388_ ( .A(\myifu/myicache/data[4][11] ), .Z(\myifu/myicache/_0498_ ) );
BUF_X1 \myifu/myicache/_3389_ ( .A(\myifu/myicache/data[5][11] ), .Z(\myifu/myicache/_0530_ ) );
BUF_X1 \myifu/myicache/_3390_ ( .A(\myifu/myicache/data[6][11] ), .Z(\myifu/myicache/_0562_ ) );
BUF_X1 \myifu/myicache/_3391_ ( .A(\myifu/myicache/data[7][11] ), .Z(\myifu/myicache/_0594_ ) );
BUF_X1 \myifu/myicache/_3392_ ( .A(\myifu/myicache/_0658_ ), .Z(\myifu/data_out [11] ) );
BUF_X1 \myifu/myicache/_3393_ ( .A(\myifu/myicache/data[0][12] ), .Z(\myifu/myicache/_0371_ ) );
BUF_X1 \myifu/myicache/_3394_ ( .A(\myifu/myicache/data[1][12] ), .Z(\myifu/myicache/_0403_ ) );
BUF_X1 \myifu/myicache/_3395_ ( .A(\myifu/myicache/data[2][12] ), .Z(\myifu/myicache/_0435_ ) );
BUF_X1 \myifu/myicache/_3396_ ( .A(\myifu/myicache/data[3][12] ), .Z(\myifu/myicache/_0467_ ) );
BUF_X1 \myifu/myicache/_3397_ ( .A(\myifu/myicache/data[4][12] ), .Z(\myifu/myicache/_0499_ ) );
BUF_X1 \myifu/myicache/_3398_ ( .A(\myifu/myicache/data[5][12] ), .Z(\myifu/myicache/_0531_ ) );
BUF_X1 \myifu/myicache/_3399_ ( .A(\myifu/myicache/data[6][12] ), .Z(\myifu/myicache/_0563_ ) );
BUF_X1 \myifu/myicache/_3400_ ( .A(\myifu/myicache/data[7][12] ), .Z(\myifu/myicache/_0595_ ) );
BUF_X1 \myifu/myicache/_3401_ ( .A(\myifu/myicache/_0659_ ), .Z(\myifu/data_out [12] ) );
BUF_X1 \myifu/myicache/_3402_ ( .A(\myifu/myicache/data[0][13] ), .Z(\myifu/myicache/_0372_ ) );
BUF_X1 \myifu/myicache/_3403_ ( .A(\myifu/myicache/data[1][13] ), .Z(\myifu/myicache/_0404_ ) );
BUF_X1 \myifu/myicache/_3404_ ( .A(\myifu/myicache/data[2][13] ), .Z(\myifu/myicache/_0436_ ) );
BUF_X1 \myifu/myicache/_3405_ ( .A(\myifu/myicache/data[3][13] ), .Z(\myifu/myicache/_0468_ ) );
BUF_X1 \myifu/myicache/_3406_ ( .A(\myifu/myicache/data[4][13] ), .Z(\myifu/myicache/_0500_ ) );
BUF_X1 \myifu/myicache/_3407_ ( .A(\myifu/myicache/data[5][13] ), .Z(\myifu/myicache/_0532_ ) );
BUF_X1 \myifu/myicache/_3408_ ( .A(\myifu/myicache/data[6][13] ), .Z(\myifu/myicache/_0564_ ) );
BUF_X1 \myifu/myicache/_3409_ ( .A(\myifu/myicache/data[7][13] ), .Z(\myifu/myicache/_0596_ ) );
BUF_X1 \myifu/myicache/_3410_ ( .A(\myifu/myicache/_0660_ ), .Z(\myifu/data_out [13] ) );
BUF_X1 \myifu/myicache/_3411_ ( .A(\myifu/myicache/data[0][14] ), .Z(\myifu/myicache/_0373_ ) );
BUF_X1 \myifu/myicache/_3412_ ( .A(\myifu/myicache/data[1][14] ), .Z(\myifu/myicache/_0405_ ) );
BUF_X1 \myifu/myicache/_3413_ ( .A(\myifu/myicache/data[2][14] ), .Z(\myifu/myicache/_0437_ ) );
BUF_X1 \myifu/myicache/_3414_ ( .A(\myifu/myicache/data[3][14] ), .Z(\myifu/myicache/_0469_ ) );
BUF_X1 \myifu/myicache/_3415_ ( .A(\myifu/myicache/data[4][14] ), .Z(\myifu/myicache/_0501_ ) );
BUF_X1 \myifu/myicache/_3416_ ( .A(\myifu/myicache/data[5][14] ), .Z(\myifu/myicache/_0533_ ) );
BUF_X1 \myifu/myicache/_3417_ ( .A(\myifu/myicache/data[6][14] ), .Z(\myifu/myicache/_0565_ ) );
BUF_X1 \myifu/myicache/_3418_ ( .A(\myifu/myicache/data[7][14] ), .Z(\myifu/myicache/_0597_ ) );
BUF_X1 \myifu/myicache/_3419_ ( .A(\myifu/myicache/_0661_ ), .Z(\myifu/data_out [14] ) );
BUF_X1 \myifu/myicache/_3420_ ( .A(\myifu/myicache/data[0][15] ), .Z(\myifu/myicache/_0374_ ) );
BUF_X1 \myifu/myicache/_3421_ ( .A(\myifu/myicache/data[1][15] ), .Z(\myifu/myicache/_0406_ ) );
BUF_X1 \myifu/myicache/_3422_ ( .A(\myifu/myicache/data[2][15] ), .Z(\myifu/myicache/_0438_ ) );
BUF_X1 \myifu/myicache/_3423_ ( .A(\myifu/myicache/data[3][15] ), .Z(\myifu/myicache/_0470_ ) );
BUF_X1 \myifu/myicache/_3424_ ( .A(\myifu/myicache/data[4][15] ), .Z(\myifu/myicache/_0502_ ) );
BUF_X1 \myifu/myicache/_3425_ ( .A(\myifu/myicache/data[5][15] ), .Z(\myifu/myicache/_0534_ ) );
BUF_X1 \myifu/myicache/_3426_ ( .A(\myifu/myicache/data[6][15] ), .Z(\myifu/myicache/_0566_ ) );
BUF_X1 \myifu/myicache/_3427_ ( .A(\myifu/myicache/data[7][15] ), .Z(\myifu/myicache/_0598_ ) );
BUF_X1 \myifu/myicache/_3428_ ( .A(\myifu/myicache/_0662_ ), .Z(\myifu/data_out [15] ) );
BUF_X1 \myifu/myicache/_3429_ ( .A(\myifu/myicache/data[0][16] ), .Z(\myifu/myicache/_0375_ ) );
BUF_X1 \myifu/myicache/_3430_ ( .A(\myifu/myicache/data[1][16] ), .Z(\myifu/myicache/_0407_ ) );
BUF_X1 \myifu/myicache/_3431_ ( .A(\myifu/myicache/data[2][16] ), .Z(\myifu/myicache/_0439_ ) );
BUF_X1 \myifu/myicache/_3432_ ( .A(\myifu/myicache/data[3][16] ), .Z(\myifu/myicache/_0471_ ) );
BUF_X1 \myifu/myicache/_3433_ ( .A(\myifu/myicache/data[4][16] ), .Z(\myifu/myicache/_0503_ ) );
BUF_X1 \myifu/myicache/_3434_ ( .A(\myifu/myicache/data[5][16] ), .Z(\myifu/myicache/_0535_ ) );
BUF_X1 \myifu/myicache/_3435_ ( .A(\myifu/myicache/data[6][16] ), .Z(\myifu/myicache/_0567_ ) );
BUF_X1 \myifu/myicache/_3436_ ( .A(\myifu/myicache/data[7][16] ), .Z(\myifu/myicache/_0599_ ) );
BUF_X1 \myifu/myicache/_3437_ ( .A(\myifu/myicache/_0663_ ), .Z(\myifu/data_out [16] ) );
BUF_X1 \myifu/myicache/_3438_ ( .A(\myifu/myicache/data[0][17] ), .Z(\myifu/myicache/_0376_ ) );
BUF_X1 \myifu/myicache/_3439_ ( .A(\myifu/myicache/data[1][17] ), .Z(\myifu/myicache/_0408_ ) );
BUF_X1 \myifu/myicache/_3440_ ( .A(\myifu/myicache/data[2][17] ), .Z(\myifu/myicache/_0440_ ) );
BUF_X1 \myifu/myicache/_3441_ ( .A(\myifu/myicache/data[3][17] ), .Z(\myifu/myicache/_0472_ ) );
BUF_X1 \myifu/myicache/_3442_ ( .A(\myifu/myicache/data[4][17] ), .Z(\myifu/myicache/_0504_ ) );
BUF_X1 \myifu/myicache/_3443_ ( .A(\myifu/myicache/data[5][17] ), .Z(\myifu/myicache/_0536_ ) );
BUF_X1 \myifu/myicache/_3444_ ( .A(\myifu/myicache/data[6][17] ), .Z(\myifu/myicache/_0568_ ) );
BUF_X1 \myifu/myicache/_3445_ ( .A(\myifu/myicache/data[7][17] ), .Z(\myifu/myicache/_0600_ ) );
BUF_X1 \myifu/myicache/_3446_ ( .A(\myifu/myicache/_0664_ ), .Z(\myifu/data_out [17] ) );
BUF_X1 \myifu/myicache/_3447_ ( .A(\myifu/myicache/data[0][18] ), .Z(\myifu/myicache/_0377_ ) );
BUF_X1 \myifu/myicache/_3448_ ( .A(\myifu/myicache/data[1][18] ), .Z(\myifu/myicache/_0409_ ) );
BUF_X1 \myifu/myicache/_3449_ ( .A(\myifu/myicache/data[2][18] ), .Z(\myifu/myicache/_0441_ ) );
BUF_X1 \myifu/myicache/_3450_ ( .A(\myifu/myicache/data[3][18] ), .Z(\myifu/myicache/_0473_ ) );
BUF_X1 \myifu/myicache/_3451_ ( .A(\myifu/myicache/data[4][18] ), .Z(\myifu/myicache/_0505_ ) );
BUF_X1 \myifu/myicache/_3452_ ( .A(\myifu/myicache/data[5][18] ), .Z(\myifu/myicache/_0537_ ) );
BUF_X1 \myifu/myicache/_3453_ ( .A(\myifu/myicache/data[6][18] ), .Z(\myifu/myicache/_0569_ ) );
BUF_X1 \myifu/myicache/_3454_ ( .A(\myifu/myicache/data[7][18] ), .Z(\myifu/myicache/_0601_ ) );
BUF_X1 \myifu/myicache/_3455_ ( .A(\myifu/myicache/_0665_ ), .Z(\myifu/data_out [18] ) );
BUF_X1 \myifu/myicache/_3456_ ( .A(\myifu/myicache/data[0][19] ), .Z(\myifu/myicache/_0378_ ) );
BUF_X1 \myifu/myicache/_3457_ ( .A(\myifu/myicache/data[1][19] ), .Z(\myifu/myicache/_0410_ ) );
BUF_X1 \myifu/myicache/_3458_ ( .A(\myifu/myicache/data[2][19] ), .Z(\myifu/myicache/_0442_ ) );
BUF_X1 \myifu/myicache/_3459_ ( .A(\myifu/myicache/data[3][19] ), .Z(\myifu/myicache/_0474_ ) );
BUF_X1 \myifu/myicache/_3460_ ( .A(\myifu/myicache/data[4][19] ), .Z(\myifu/myicache/_0506_ ) );
BUF_X1 \myifu/myicache/_3461_ ( .A(\myifu/myicache/data[5][19] ), .Z(\myifu/myicache/_0538_ ) );
BUF_X1 \myifu/myicache/_3462_ ( .A(\myifu/myicache/data[6][19] ), .Z(\myifu/myicache/_0570_ ) );
BUF_X1 \myifu/myicache/_3463_ ( .A(\myifu/myicache/data[7][19] ), .Z(\myifu/myicache/_0602_ ) );
BUF_X1 \myifu/myicache/_3464_ ( .A(\myifu/myicache/_0666_ ), .Z(\myifu/data_out [19] ) );
BUF_X1 \myifu/myicache/_3465_ ( .A(\myifu/myicache/data[0][20] ), .Z(\myifu/myicache/_0380_ ) );
BUF_X1 \myifu/myicache/_3466_ ( .A(\myifu/myicache/data[1][20] ), .Z(\myifu/myicache/_0412_ ) );
BUF_X1 \myifu/myicache/_3467_ ( .A(\myifu/myicache/data[2][20] ), .Z(\myifu/myicache/_0444_ ) );
BUF_X1 \myifu/myicache/_3468_ ( .A(\myifu/myicache/data[3][20] ), .Z(\myifu/myicache/_0476_ ) );
BUF_X1 \myifu/myicache/_3469_ ( .A(\myifu/myicache/data[4][20] ), .Z(\myifu/myicache/_0508_ ) );
BUF_X1 \myifu/myicache/_3470_ ( .A(\myifu/myicache/data[5][20] ), .Z(\myifu/myicache/_0540_ ) );
BUF_X1 \myifu/myicache/_3471_ ( .A(\myifu/myicache/data[6][20] ), .Z(\myifu/myicache/_0572_ ) );
BUF_X1 \myifu/myicache/_3472_ ( .A(\myifu/myicache/data[7][20] ), .Z(\myifu/myicache/_0604_ ) );
BUF_X1 \myifu/myicache/_3473_ ( .A(\myifu/myicache/_0668_ ), .Z(\myifu/data_out [20] ) );
BUF_X1 \myifu/myicache/_3474_ ( .A(\myifu/myicache/data[0][21] ), .Z(\myifu/myicache/_0381_ ) );
BUF_X1 \myifu/myicache/_3475_ ( .A(\myifu/myicache/data[1][21] ), .Z(\myifu/myicache/_0413_ ) );
BUF_X1 \myifu/myicache/_3476_ ( .A(\myifu/myicache/data[2][21] ), .Z(\myifu/myicache/_0445_ ) );
BUF_X1 \myifu/myicache/_3477_ ( .A(\myifu/myicache/data[3][21] ), .Z(\myifu/myicache/_0477_ ) );
BUF_X1 \myifu/myicache/_3478_ ( .A(\myifu/myicache/data[4][21] ), .Z(\myifu/myicache/_0509_ ) );
BUF_X1 \myifu/myicache/_3479_ ( .A(\myifu/myicache/data[5][21] ), .Z(\myifu/myicache/_0541_ ) );
BUF_X1 \myifu/myicache/_3480_ ( .A(\myifu/myicache/data[6][21] ), .Z(\myifu/myicache/_0573_ ) );
BUF_X1 \myifu/myicache/_3481_ ( .A(\myifu/myicache/data[7][21] ), .Z(\myifu/myicache/_0605_ ) );
BUF_X1 \myifu/myicache/_3482_ ( .A(\myifu/myicache/_0669_ ), .Z(\myifu/data_out [21] ) );
BUF_X1 \myifu/myicache/_3483_ ( .A(\myifu/myicache/data[0][22] ), .Z(\myifu/myicache/_0382_ ) );
BUF_X1 \myifu/myicache/_3484_ ( .A(\myifu/myicache/data[1][22] ), .Z(\myifu/myicache/_0414_ ) );
BUF_X1 \myifu/myicache/_3485_ ( .A(\myifu/myicache/data[2][22] ), .Z(\myifu/myicache/_0446_ ) );
BUF_X1 \myifu/myicache/_3486_ ( .A(\myifu/myicache/data[3][22] ), .Z(\myifu/myicache/_0478_ ) );
BUF_X1 \myifu/myicache/_3487_ ( .A(\myifu/myicache/data[4][22] ), .Z(\myifu/myicache/_0510_ ) );
BUF_X1 \myifu/myicache/_3488_ ( .A(\myifu/myicache/data[5][22] ), .Z(\myifu/myicache/_0542_ ) );
BUF_X1 \myifu/myicache/_3489_ ( .A(\myifu/myicache/data[6][22] ), .Z(\myifu/myicache/_0574_ ) );
BUF_X1 \myifu/myicache/_3490_ ( .A(\myifu/myicache/data[7][22] ), .Z(\myifu/myicache/_0606_ ) );
BUF_X1 \myifu/myicache/_3491_ ( .A(\myifu/myicache/_0670_ ), .Z(\myifu/data_out [22] ) );
BUF_X1 \myifu/myicache/_3492_ ( .A(\myifu/myicache/data[0][23] ), .Z(\myifu/myicache/_0383_ ) );
BUF_X1 \myifu/myicache/_3493_ ( .A(\myifu/myicache/data[1][23] ), .Z(\myifu/myicache/_0415_ ) );
BUF_X1 \myifu/myicache/_3494_ ( .A(\myifu/myicache/data[2][23] ), .Z(\myifu/myicache/_0447_ ) );
BUF_X1 \myifu/myicache/_3495_ ( .A(\myifu/myicache/data[3][23] ), .Z(\myifu/myicache/_0479_ ) );
BUF_X1 \myifu/myicache/_3496_ ( .A(\myifu/myicache/data[4][23] ), .Z(\myifu/myicache/_0511_ ) );
BUF_X1 \myifu/myicache/_3497_ ( .A(\myifu/myicache/data[5][23] ), .Z(\myifu/myicache/_0543_ ) );
BUF_X1 \myifu/myicache/_3498_ ( .A(\myifu/myicache/data[6][23] ), .Z(\myifu/myicache/_0575_ ) );
BUF_X1 \myifu/myicache/_3499_ ( .A(\myifu/myicache/data[7][23] ), .Z(\myifu/myicache/_0607_ ) );
BUF_X1 \myifu/myicache/_3500_ ( .A(\myifu/myicache/_0671_ ), .Z(\myifu/data_out [23] ) );
BUF_X1 \myifu/myicache/_3501_ ( .A(\myifu/myicache/data[0][24] ), .Z(\myifu/myicache/_0384_ ) );
BUF_X1 \myifu/myicache/_3502_ ( .A(\myifu/myicache/data[1][24] ), .Z(\myifu/myicache/_0416_ ) );
BUF_X1 \myifu/myicache/_3503_ ( .A(\myifu/myicache/data[2][24] ), .Z(\myifu/myicache/_0448_ ) );
BUF_X1 \myifu/myicache/_3504_ ( .A(\myifu/myicache/data[3][24] ), .Z(\myifu/myicache/_0480_ ) );
BUF_X1 \myifu/myicache/_3505_ ( .A(\myifu/myicache/data[4][24] ), .Z(\myifu/myicache/_0512_ ) );
BUF_X1 \myifu/myicache/_3506_ ( .A(\myifu/myicache/data[5][24] ), .Z(\myifu/myicache/_0544_ ) );
BUF_X1 \myifu/myicache/_3507_ ( .A(\myifu/myicache/data[6][24] ), .Z(\myifu/myicache/_0576_ ) );
BUF_X1 \myifu/myicache/_3508_ ( .A(\myifu/myicache/data[7][24] ), .Z(\myifu/myicache/_0608_ ) );
BUF_X1 \myifu/myicache/_3509_ ( .A(\myifu/myicache/_0672_ ), .Z(\myifu/data_out [24] ) );
BUF_X1 \myifu/myicache/_3510_ ( .A(\myifu/myicache/data[0][25] ), .Z(\myifu/myicache/_0385_ ) );
BUF_X1 \myifu/myicache/_3511_ ( .A(\myifu/myicache/data[1][25] ), .Z(\myifu/myicache/_0417_ ) );
BUF_X1 \myifu/myicache/_3512_ ( .A(\myifu/myicache/data[2][25] ), .Z(\myifu/myicache/_0449_ ) );
BUF_X1 \myifu/myicache/_3513_ ( .A(\myifu/myicache/data[3][25] ), .Z(\myifu/myicache/_0481_ ) );
BUF_X1 \myifu/myicache/_3514_ ( .A(\myifu/myicache/data[4][25] ), .Z(\myifu/myicache/_0513_ ) );
BUF_X1 \myifu/myicache/_3515_ ( .A(\myifu/myicache/data[5][25] ), .Z(\myifu/myicache/_0545_ ) );
BUF_X1 \myifu/myicache/_3516_ ( .A(\myifu/myicache/data[6][25] ), .Z(\myifu/myicache/_0577_ ) );
BUF_X1 \myifu/myicache/_3517_ ( .A(\myifu/myicache/data[7][25] ), .Z(\myifu/myicache/_0609_ ) );
BUF_X1 \myifu/myicache/_3518_ ( .A(\myifu/myicache/_0673_ ), .Z(\myifu/data_out [25] ) );
BUF_X1 \myifu/myicache/_3519_ ( .A(\myifu/myicache/data[0][26] ), .Z(\myifu/myicache/_0386_ ) );
BUF_X1 \myifu/myicache/_3520_ ( .A(\myifu/myicache/data[1][26] ), .Z(\myifu/myicache/_0418_ ) );
BUF_X1 \myifu/myicache/_3521_ ( .A(\myifu/myicache/data[2][26] ), .Z(\myifu/myicache/_0450_ ) );
BUF_X1 \myifu/myicache/_3522_ ( .A(\myifu/myicache/data[3][26] ), .Z(\myifu/myicache/_0482_ ) );
BUF_X1 \myifu/myicache/_3523_ ( .A(\myifu/myicache/data[4][26] ), .Z(\myifu/myicache/_0514_ ) );
BUF_X1 \myifu/myicache/_3524_ ( .A(\myifu/myicache/data[5][26] ), .Z(\myifu/myicache/_0546_ ) );
BUF_X1 \myifu/myicache/_3525_ ( .A(\myifu/myicache/data[6][26] ), .Z(\myifu/myicache/_0578_ ) );
BUF_X1 \myifu/myicache/_3526_ ( .A(\myifu/myicache/data[7][26] ), .Z(\myifu/myicache/_0610_ ) );
BUF_X1 \myifu/myicache/_3527_ ( .A(\myifu/myicache/_0674_ ), .Z(\myifu/data_out [26] ) );
BUF_X1 \myifu/myicache/_3528_ ( .A(\myifu/myicache/data[0][27] ), .Z(\myifu/myicache/_0387_ ) );
BUF_X1 \myifu/myicache/_3529_ ( .A(\myifu/myicache/data[1][27] ), .Z(\myifu/myicache/_0419_ ) );
BUF_X1 \myifu/myicache/_3530_ ( .A(\myifu/myicache/data[2][27] ), .Z(\myifu/myicache/_0451_ ) );
BUF_X1 \myifu/myicache/_3531_ ( .A(\myifu/myicache/data[3][27] ), .Z(\myifu/myicache/_0483_ ) );
BUF_X1 \myifu/myicache/_3532_ ( .A(\myifu/myicache/data[4][27] ), .Z(\myifu/myicache/_0515_ ) );
BUF_X1 \myifu/myicache/_3533_ ( .A(\myifu/myicache/data[5][27] ), .Z(\myifu/myicache/_0547_ ) );
BUF_X1 \myifu/myicache/_3534_ ( .A(\myifu/myicache/data[6][27] ), .Z(\myifu/myicache/_0579_ ) );
BUF_X1 \myifu/myicache/_3535_ ( .A(\myifu/myicache/data[7][27] ), .Z(\myifu/myicache/_0611_ ) );
BUF_X1 \myifu/myicache/_3536_ ( .A(\myifu/myicache/_0675_ ), .Z(\myifu/data_out [27] ) );
BUF_X1 \myifu/myicache/_3537_ ( .A(\myifu/myicache/data[0][28] ), .Z(\myifu/myicache/_0388_ ) );
BUF_X1 \myifu/myicache/_3538_ ( .A(\myifu/myicache/data[1][28] ), .Z(\myifu/myicache/_0420_ ) );
BUF_X1 \myifu/myicache/_3539_ ( .A(\myifu/myicache/data[2][28] ), .Z(\myifu/myicache/_0452_ ) );
BUF_X1 \myifu/myicache/_3540_ ( .A(\myifu/myicache/data[3][28] ), .Z(\myifu/myicache/_0484_ ) );
BUF_X1 \myifu/myicache/_3541_ ( .A(\myifu/myicache/data[4][28] ), .Z(\myifu/myicache/_0516_ ) );
BUF_X1 \myifu/myicache/_3542_ ( .A(\myifu/myicache/data[5][28] ), .Z(\myifu/myicache/_0548_ ) );
BUF_X1 \myifu/myicache/_3543_ ( .A(\myifu/myicache/data[6][28] ), .Z(\myifu/myicache/_0580_ ) );
BUF_X1 \myifu/myicache/_3544_ ( .A(\myifu/myicache/data[7][28] ), .Z(\myifu/myicache/_0612_ ) );
BUF_X1 \myifu/myicache/_3545_ ( .A(\myifu/myicache/_0676_ ), .Z(\myifu/data_out [28] ) );
BUF_X1 \myifu/myicache/_3546_ ( .A(\myifu/myicache/data[0][29] ), .Z(\myifu/myicache/_0389_ ) );
BUF_X1 \myifu/myicache/_3547_ ( .A(\myifu/myicache/data[1][29] ), .Z(\myifu/myicache/_0421_ ) );
BUF_X1 \myifu/myicache/_3548_ ( .A(\myifu/myicache/data[2][29] ), .Z(\myifu/myicache/_0453_ ) );
BUF_X1 \myifu/myicache/_3549_ ( .A(\myifu/myicache/data[3][29] ), .Z(\myifu/myicache/_0485_ ) );
BUF_X1 \myifu/myicache/_3550_ ( .A(\myifu/myicache/data[4][29] ), .Z(\myifu/myicache/_0517_ ) );
BUF_X1 \myifu/myicache/_3551_ ( .A(\myifu/myicache/data[5][29] ), .Z(\myifu/myicache/_0549_ ) );
BUF_X1 \myifu/myicache/_3552_ ( .A(\myifu/myicache/data[6][29] ), .Z(\myifu/myicache/_0581_ ) );
BUF_X1 \myifu/myicache/_3553_ ( .A(\myifu/myicache/data[7][29] ), .Z(\myifu/myicache/_0613_ ) );
BUF_X1 \myifu/myicache/_3554_ ( .A(\myifu/myicache/_0677_ ), .Z(\myifu/data_out [29] ) );
BUF_X1 \myifu/myicache/_3555_ ( .A(\myifu/myicache/data[0][30] ), .Z(\myifu/myicache/_0391_ ) );
BUF_X1 \myifu/myicache/_3556_ ( .A(\myifu/myicache/data[1][30] ), .Z(\myifu/myicache/_0423_ ) );
BUF_X1 \myifu/myicache/_3557_ ( .A(\myifu/myicache/data[2][30] ), .Z(\myifu/myicache/_0455_ ) );
BUF_X1 \myifu/myicache/_3558_ ( .A(\myifu/myicache/data[3][30] ), .Z(\myifu/myicache/_0487_ ) );
BUF_X1 \myifu/myicache/_3559_ ( .A(\myifu/myicache/data[4][30] ), .Z(\myifu/myicache/_0519_ ) );
BUF_X1 \myifu/myicache/_3560_ ( .A(\myifu/myicache/data[5][30] ), .Z(\myifu/myicache/_0551_ ) );
BUF_X1 \myifu/myicache/_3561_ ( .A(\myifu/myicache/data[6][30] ), .Z(\myifu/myicache/_0583_ ) );
BUF_X1 \myifu/myicache/_3562_ ( .A(\myifu/myicache/data[7][30] ), .Z(\myifu/myicache/_0615_ ) );
BUF_X1 \myifu/myicache/_3563_ ( .A(\myifu/myicache/_0679_ ), .Z(\myifu/data_out [30] ) );
BUF_X1 \myifu/myicache/_3564_ ( .A(\myifu/myicache/data[0][31] ), .Z(\myifu/myicache/_0392_ ) );
BUF_X1 \myifu/myicache/_3565_ ( .A(\myifu/myicache/data[1][31] ), .Z(\myifu/myicache/_0424_ ) );
BUF_X1 \myifu/myicache/_3566_ ( .A(\myifu/myicache/data[2][31] ), .Z(\myifu/myicache/_0456_ ) );
BUF_X1 \myifu/myicache/_3567_ ( .A(\myifu/myicache/data[3][31] ), .Z(\myifu/myicache/_0488_ ) );
BUF_X1 \myifu/myicache/_3568_ ( .A(\myifu/myicache/data[4][31] ), .Z(\myifu/myicache/_0520_ ) );
BUF_X1 \myifu/myicache/_3569_ ( .A(\myifu/myicache/data[5][31] ), .Z(\myifu/myicache/_0552_ ) );
BUF_X1 \myifu/myicache/_3570_ ( .A(\myifu/myicache/data[6][31] ), .Z(\myifu/myicache/_0584_ ) );
BUF_X1 \myifu/myicache/_3571_ ( .A(\myifu/myicache/data[7][31] ), .Z(\myifu/myicache/_0616_ ) );
BUF_X1 \myifu/myicache/_3572_ ( .A(\myifu/myicache/_0680_ ), .Z(\myifu/data_out [31] ) );
BUF_X1 \myifu/myicache/_3573_ ( .A(\rdata_IFU [0] ), .Z(\myifu/myicache/_0624_ ) );
BUF_X1 \myifu/myicache/_3574_ ( .A(\myifu/myicache/_0000_ ), .Z(\myifu/myicache/_1602_ ) );
BUF_X1 \myifu/myicache/_3575_ ( .A(\rdata_IFU [1] ), .Z(\myifu/myicache/_0635_ ) );
BUF_X1 \myifu/myicache/_3576_ ( .A(\myifu/myicache/_0001_ ), .Z(\myifu/myicache/_1603_ ) );
BUF_X1 \myifu/myicache/_3577_ ( .A(\rdata_IFU [2] ), .Z(\myifu/myicache/_0646_ ) );
BUF_X1 \myifu/myicache/_3578_ ( .A(\myifu/myicache/_0002_ ), .Z(\myifu/myicache/_1604_ ) );
BUF_X1 \myifu/myicache/_3579_ ( .A(\rdata_IFU [3] ), .Z(\myifu/myicache/_0649_ ) );
BUF_X1 \myifu/myicache/_3580_ ( .A(\myifu/myicache/_0003_ ), .Z(\myifu/myicache/_1605_ ) );
BUF_X1 \myifu/myicache/_3581_ ( .A(\rdata_IFU [4] ), .Z(\myifu/myicache/_0650_ ) );
BUF_X1 \myifu/myicache/_3582_ ( .A(\myifu/myicache/_0004_ ), .Z(\myifu/myicache/_1606_ ) );
BUF_X1 \myifu/myicache/_3583_ ( .A(\rdata_IFU [5] ), .Z(\myifu/myicache/_0651_ ) );
BUF_X1 \myifu/myicache/_3584_ ( .A(\myifu/myicache/_0005_ ), .Z(\myifu/myicache/_1607_ ) );
BUF_X1 \myifu/myicache/_3585_ ( .A(\rdata_IFU [6] ), .Z(\myifu/myicache/_0652_ ) );
BUF_X1 \myifu/myicache/_3586_ ( .A(\myifu/myicache/_0006_ ), .Z(\myifu/myicache/_1608_ ) );
BUF_X1 \myifu/myicache/_3587_ ( .A(\rdata_IFU [7] ), .Z(\myifu/myicache/_0653_ ) );
BUF_X1 \myifu/myicache/_3588_ ( .A(\myifu/myicache/_0007_ ), .Z(\myifu/myicache/_1609_ ) );
BUF_X1 \myifu/myicache/_3589_ ( .A(\rdata_IFU [8] ), .Z(\myifu/myicache/_0654_ ) );
BUF_X1 \myifu/myicache/_3590_ ( .A(\myifu/myicache/_0008_ ), .Z(\myifu/myicache/_1610_ ) );
BUF_X1 \myifu/myicache/_3591_ ( .A(\rdata_IFU [9] ), .Z(\myifu/myicache/_0655_ ) );
BUF_X1 \myifu/myicache/_3592_ ( .A(\myifu/myicache/_0009_ ), .Z(\myifu/myicache/_1611_ ) );
BUF_X1 \myifu/myicache/_3593_ ( .A(\rdata_IFU [10] ), .Z(\myifu/myicache/_0625_ ) );
BUF_X1 \myifu/myicache/_3594_ ( .A(\myifu/myicache/_0010_ ), .Z(\myifu/myicache/_1612_ ) );
BUF_X1 \myifu/myicache/_3595_ ( .A(\rdata_IFU [11] ), .Z(\myifu/myicache/_0626_ ) );
BUF_X1 \myifu/myicache/_3596_ ( .A(\myifu/myicache/_0011_ ), .Z(\myifu/myicache/_1613_ ) );
BUF_X1 \myifu/myicache/_3597_ ( .A(\rdata_IFU [12] ), .Z(\myifu/myicache/_0627_ ) );
BUF_X1 \myifu/myicache/_3598_ ( .A(\myifu/myicache/_0012_ ), .Z(\myifu/myicache/_1614_ ) );
BUF_X1 \myifu/myicache/_3599_ ( .A(\rdata_IFU [13] ), .Z(\myifu/myicache/_0628_ ) );
BUF_X1 \myifu/myicache/_3600_ ( .A(\myifu/myicache/_0013_ ), .Z(\myifu/myicache/_1615_ ) );
BUF_X1 \myifu/myicache/_3601_ ( .A(\rdata_IFU [14] ), .Z(\myifu/myicache/_0629_ ) );
BUF_X1 \myifu/myicache/_3602_ ( .A(\myifu/myicache/_0014_ ), .Z(\myifu/myicache/_1616_ ) );
BUF_X1 \myifu/myicache/_3603_ ( .A(\rdata_IFU [15] ), .Z(\myifu/myicache/_0630_ ) );
BUF_X1 \myifu/myicache/_3604_ ( .A(\myifu/myicache/_0015_ ), .Z(\myifu/myicache/_1617_ ) );
BUF_X1 \myifu/myicache/_3605_ ( .A(\rdata_IFU [16] ), .Z(\myifu/myicache/_0631_ ) );
BUF_X1 \myifu/myicache/_3606_ ( .A(\myifu/myicache/_0016_ ), .Z(\myifu/myicache/_1618_ ) );
BUF_X1 \myifu/myicache/_3607_ ( .A(\rdata_IFU [17] ), .Z(\myifu/myicache/_0632_ ) );
BUF_X1 \myifu/myicache/_3608_ ( .A(\myifu/myicache/_0017_ ), .Z(\myifu/myicache/_1619_ ) );
BUF_X1 \myifu/myicache/_3609_ ( .A(\rdata_IFU [18] ), .Z(\myifu/myicache/_0633_ ) );
BUF_X1 \myifu/myicache/_3610_ ( .A(\myifu/myicache/_0018_ ), .Z(\myifu/myicache/_1620_ ) );
BUF_X1 \myifu/myicache/_3611_ ( .A(\rdata_IFU [19] ), .Z(\myifu/myicache/_0634_ ) );
BUF_X1 \myifu/myicache/_3612_ ( .A(\myifu/myicache/_0019_ ), .Z(\myifu/myicache/_1621_ ) );
BUF_X1 \myifu/myicache/_3613_ ( .A(\rdata_IFU [20] ), .Z(\myifu/myicache/_0636_ ) );
BUF_X1 \myifu/myicache/_3614_ ( .A(\myifu/myicache/_0020_ ), .Z(\myifu/myicache/_1622_ ) );
BUF_X1 \myifu/myicache/_3615_ ( .A(\rdata_IFU [21] ), .Z(\myifu/myicache/_0637_ ) );
BUF_X1 \myifu/myicache/_3616_ ( .A(\myifu/myicache/_0021_ ), .Z(\myifu/myicache/_1623_ ) );
BUF_X1 \myifu/myicache/_3617_ ( .A(\rdata_IFU [22] ), .Z(\myifu/myicache/_0638_ ) );
BUF_X1 \myifu/myicache/_3618_ ( .A(\myifu/myicache/_0022_ ), .Z(\myifu/myicache/_1624_ ) );
BUF_X1 \myifu/myicache/_3619_ ( .A(\rdata_IFU [23] ), .Z(\myifu/myicache/_0639_ ) );
BUF_X1 \myifu/myicache/_3620_ ( .A(\myifu/myicache/_0023_ ), .Z(\myifu/myicache/_1625_ ) );
BUF_X1 \myifu/myicache/_3621_ ( .A(\rdata_IFU [24] ), .Z(\myifu/myicache/_0640_ ) );
BUF_X1 \myifu/myicache/_3622_ ( .A(\myifu/myicache/_0024_ ), .Z(\myifu/myicache/_1626_ ) );
BUF_X1 \myifu/myicache/_3623_ ( .A(\rdata_IFU [25] ), .Z(\myifu/myicache/_0641_ ) );
BUF_X1 \myifu/myicache/_3624_ ( .A(\myifu/myicache/_0025_ ), .Z(\myifu/myicache/_1627_ ) );
BUF_X1 \myifu/myicache/_3625_ ( .A(\rdata_IFU [26] ), .Z(\myifu/myicache/_0642_ ) );
BUF_X1 \myifu/myicache/_3626_ ( .A(\myifu/myicache/_0026_ ), .Z(\myifu/myicache/_1628_ ) );
BUF_X1 \myifu/myicache/_3627_ ( .A(\rdata_IFU [27] ), .Z(\myifu/myicache/_0643_ ) );
BUF_X1 \myifu/myicache/_3628_ ( .A(\myifu/myicache/_0027_ ), .Z(\myifu/myicache/_1629_ ) );
BUF_X1 \myifu/myicache/_3629_ ( .A(\rdata_IFU [28] ), .Z(\myifu/myicache/_0644_ ) );
BUF_X1 \myifu/myicache/_3630_ ( .A(\myifu/myicache/_0028_ ), .Z(\myifu/myicache/_1630_ ) );
BUF_X1 \myifu/myicache/_3631_ ( .A(\rdata_IFU [29] ), .Z(\myifu/myicache/_0645_ ) );
BUF_X1 \myifu/myicache/_3632_ ( .A(\myifu/myicache/_0029_ ), .Z(\myifu/myicache/_1631_ ) );
BUF_X1 \myifu/myicache/_3633_ ( .A(\rdata_IFU [30] ), .Z(\myifu/myicache/_0647_ ) );
BUF_X1 \myifu/myicache/_3634_ ( .A(\myifu/myicache/_0030_ ), .Z(\myifu/myicache/_1632_ ) );
BUF_X1 \myifu/myicache/_3635_ ( .A(\rdata_IFU [31] ), .Z(\myifu/myicache/_0648_ ) );
BUF_X1 \myifu/myicache/_3636_ ( .A(\myifu/myicache/_0031_ ), .Z(\myifu/myicache/_1633_ ) );
BUF_X1 \myifu/myicache/_3637_ ( .A(\myifu/myicache/_0032_ ), .Z(\myifu/myicache/_1634_ ) );
BUF_X1 \myifu/myicache/_3638_ ( .A(\myifu/myicache/_0033_ ), .Z(\myifu/myicache/_1635_ ) );
BUF_X1 \myifu/myicache/_3639_ ( .A(\myifu/myicache/_0034_ ), .Z(\myifu/myicache/_1636_ ) );
BUF_X1 \myifu/myicache/_3640_ ( .A(\myifu/myicache/_0035_ ), .Z(\myifu/myicache/_1637_ ) );
BUF_X1 \myifu/myicache/_3641_ ( .A(\myifu/myicache/_0036_ ), .Z(\myifu/myicache/_1638_ ) );
BUF_X1 \myifu/myicache/_3642_ ( .A(\myifu/myicache/_0037_ ), .Z(\myifu/myicache/_1639_ ) );
BUF_X1 \myifu/myicache/_3643_ ( .A(\myifu/myicache/_0038_ ), .Z(\myifu/myicache/_1640_ ) );
BUF_X1 \myifu/myicache/_3644_ ( .A(\myifu/myicache/_0039_ ), .Z(\myifu/myicache/_1641_ ) );
BUF_X1 \myifu/myicache/_3645_ ( .A(\myifu/myicache/_0040_ ), .Z(\myifu/myicache/_1642_ ) );
BUF_X1 \myifu/myicache/_3646_ ( .A(\myifu/myicache/_0041_ ), .Z(\myifu/myicache/_1643_ ) );
BUF_X1 \myifu/myicache/_3647_ ( .A(\myifu/myicache/_0042_ ), .Z(\myifu/myicache/_1644_ ) );
BUF_X1 \myifu/myicache/_3648_ ( .A(\myifu/myicache/_0043_ ), .Z(\myifu/myicache/_1645_ ) );
BUF_X1 \myifu/myicache/_3649_ ( .A(\myifu/myicache/_0044_ ), .Z(\myifu/myicache/_1646_ ) );
BUF_X1 \myifu/myicache/_3650_ ( .A(\myifu/myicache/_0045_ ), .Z(\myifu/myicache/_1647_ ) );
BUF_X1 \myifu/myicache/_3651_ ( .A(\myifu/myicache/_0046_ ), .Z(\myifu/myicache/_1648_ ) );
BUF_X1 \myifu/myicache/_3652_ ( .A(\myifu/myicache/_0047_ ), .Z(\myifu/myicache/_1649_ ) );
BUF_X1 \myifu/myicache/_3653_ ( .A(\myifu/myicache/_0048_ ), .Z(\myifu/myicache/_1650_ ) );
BUF_X1 \myifu/myicache/_3654_ ( .A(\myifu/myicache/_0049_ ), .Z(\myifu/myicache/_1651_ ) );
BUF_X1 \myifu/myicache/_3655_ ( .A(\myifu/myicache/_0050_ ), .Z(\myifu/myicache/_1652_ ) );
BUF_X1 \myifu/myicache/_3656_ ( .A(\myifu/myicache/_0051_ ), .Z(\myifu/myicache/_1653_ ) );
BUF_X1 \myifu/myicache/_3657_ ( .A(\myifu/myicache/_0052_ ), .Z(\myifu/myicache/_1654_ ) );
BUF_X1 \myifu/myicache/_3658_ ( .A(\myifu/myicache/_0053_ ), .Z(\myifu/myicache/_1655_ ) );
BUF_X1 \myifu/myicache/_3659_ ( .A(\myifu/myicache/_0054_ ), .Z(\myifu/myicache/_1656_ ) );
BUF_X1 \myifu/myicache/_3660_ ( .A(\myifu/myicache/_0055_ ), .Z(\myifu/myicache/_1657_ ) );
BUF_X1 \myifu/myicache/_3661_ ( .A(\myifu/myicache/_0056_ ), .Z(\myifu/myicache/_1658_ ) );
BUF_X1 \myifu/myicache/_3662_ ( .A(\myifu/myicache/_0057_ ), .Z(\myifu/myicache/_1659_ ) );
BUF_X1 \myifu/myicache/_3663_ ( .A(\myifu/myicache/_0058_ ), .Z(\myifu/myicache/_1660_ ) );
BUF_X1 \myifu/myicache/_3664_ ( .A(\myifu/myicache/_0059_ ), .Z(\myifu/myicache/_1661_ ) );
BUF_X1 \myifu/myicache/_3665_ ( .A(\myifu/myicache/_0060_ ), .Z(\myifu/myicache/_1662_ ) );
BUF_X1 \myifu/myicache/_3666_ ( .A(\myifu/myicache/_0061_ ), .Z(\myifu/myicache/_1663_ ) );
BUF_X1 \myifu/myicache/_3667_ ( .A(\myifu/myicache/_0062_ ), .Z(\myifu/myicache/_1664_ ) );
BUF_X1 \myifu/myicache/_3668_ ( .A(\myifu/myicache/_0063_ ), .Z(\myifu/myicache/_1665_ ) );
BUF_X1 \myifu/myicache/_3669_ ( .A(\myifu/myicache/_0064_ ), .Z(\myifu/myicache/_1666_ ) );
BUF_X1 \myifu/myicache/_3670_ ( .A(\myifu/myicache/_0065_ ), .Z(\myifu/myicache/_1667_ ) );
BUF_X1 \myifu/myicache/_3671_ ( .A(\myifu/myicache/_0066_ ), .Z(\myifu/myicache/_1668_ ) );
BUF_X1 \myifu/myicache/_3672_ ( .A(\myifu/myicache/_0067_ ), .Z(\myifu/myicache/_1669_ ) );
BUF_X1 \myifu/myicache/_3673_ ( .A(\myifu/myicache/_0068_ ), .Z(\myifu/myicache/_1670_ ) );
BUF_X1 \myifu/myicache/_3674_ ( .A(\myifu/myicache/_0069_ ), .Z(\myifu/myicache/_1671_ ) );
BUF_X1 \myifu/myicache/_3675_ ( .A(\myifu/myicache/_0070_ ), .Z(\myifu/myicache/_1672_ ) );
BUF_X1 \myifu/myicache/_3676_ ( .A(\myifu/myicache/_0071_ ), .Z(\myifu/myicache/_1673_ ) );
BUF_X1 \myifu/myicache/_3677_ ( .A(\myifu/myicache/_0072_ ), .Z(\myifu/myicache/_1674_ ) );
BUF_X1 \myifu/myicache/_3678_ ( .A(\myifu/myicache/_0073_ ), .Z(\myifu/myicache/_1675_ ) );
BUF_X1 \myifu/myicache/_3679_ ( .A(\myifu/myicache/_0074_ ), .Z(\myifu/myicache/_1676_ ) );
BUF_X1 \myifu/myicache/_3680_ ( .A(\myifu/myicache/_0075_ ), .Z(\myifu/myicache/_1677_ ) );
BUF_X1 \myifu/myicache/_3681_ ( .A(\myifu/myicache/_0076_ ), .Z(\myifu/myicache/_1678_ ) );
BUF_X1 \myifu/myicache/_3682_ ( .A(\myifu/myicache/_0077_ ), .Z(\myifu/myicache/_1679_ ) );
BUF_X1 \myifu/myicache/_3683_ ( .A(\myifu/myicache/_0078_ ), .Z(\myifu/myicache/_1680_ ) );
BUF_X1 \myifu/myicache/_3684_ ( .A(\myifu/myicache/_0079_ ), .Z(\myifu/myicache/_1681_ ) );
BUF_X1 \myifu/myicache/_3685_ ( .A(\myifu/myicache/_0080_ ), .Z(\myifu/myicache/_1682_ ) );
BUF_X1 \myifu/myicache/_3686_ ( .A(\myifu/myicache/_0081_ ), .Z(\myifu/myicache/_1683_ ) );
BUF_X1 \myifu/myicache/_3687_ ( .A(\myifu/myicache/_0082_ ), .Z(\myifu/myicache/_1684_ ) );
BUF_X1 \myifu/myicache/_3688_ ( .A(\myifu/myicache/_0083_ ), .Z(\myifu/myicache/_1685_ ) );
BUF_X1 \myifu/myicache/_3689_ ( .A(\myifu/myicache/_0084_ ), .Z(\myifu/myicache/_1686_ ) );
BUF_X1 \myifu/myicache/_3690_ ( .A(\myifu/myicache/_0085_ ), .Z(\myifu/myicache/_1687_ ) );
BUF_X1 \myifu/myicache/_3691_ ( .A(\myifu/myicache/_0086_ ), .Z(\myifu/myicache/_1688_ ) );
BUF_X1 \myifu/myicache/_3692_ ( .A(\myifu/myicache/_0087_ ), .Z(\myifu/myicache/_1689_ ) );
BUF_X1 \myifu/myicache/_3693_ ( .A(\myifu/myicache/_0088_ ), .Z(\myifu/myicache/_1690_ ) );
BUF_X1 \myifu/myicache/_3694_ ( .A(\myifu/myicache/_0089_ ), .Z(\myifu/myicache/_1691_ ) );
BUF_X1 \myifu/myicache/_3695_ ( .A(\myifu/myicache/_0090_ ), .Z(\myifu/myicache/_1692_ ) );
BUF_X1 \myifu/myicache/_3696_ ( .A(\myifu/myicache/_0091_ ), .Z(\myifu/myicache/_1693_ ) );
BUF_X1 \myifu/myicache/_3697_ ( .A(\myifu/myicache/_0092_ ), .Z(\myifu/myicache/_1694_ ) );
BUF_X1 \myifu/myicache/_3698_ ( .A(\myifu/myicache/_0093_ ), .Z(\myifu/myicache/_1695_ ) );
BUF_X1 \myifu/myicache/_3699_ ( .A(\myifu/myicache/_0094_ ), .Z(\myifu/myicache/_1696_ ) );
BUF_X1 \myifu/myicache/_3700_ ( .A(\myifu/myicache/_0095_ ), .Z(\myifu/myicache/_1697_ ) );
BUF_X1 \myifu/myicache/_3701_ ( .A(\myifu/myicache/_0096_ ), .Z(\myifu/myicache/_1698_ ) );
BUF_X1 \myifu/myicache/_3702_ ( .A(\myifu/myicache/_0097_ ), .Z(\myifu/myicache/_1699_ ) );
BUF_X1 \myifu/myicache/_3703_ ( .A(\myifu/myicache/_0098_ ), .Z(\myifu/myicache/_1700_ ) );
BUF_X1 \myifu/myicache/_3704_ ( .A(\myifu/myicache/_0099_ ), .Z(\myifu/myicache/_1701_ ) );
BUF_X1 \myifu/myicache/_3705_ ( .A(\myifu/myicache/_0100_ ), .Z(\myifu/myicache/_1702_ ) );
BUF_X1 \myifu/myicache/_3706_ ( .A(\myifu/myicache/_0101_ ), .Z(\myifu/myicache/_1703_ ) );
BUF_X1 \myifu/myicache/_3707_ ( .A(\myifu/myicache/_0102_ ), .Z(\myifu/myicache/_1704_ ) );
BUF_X1 \myifu/myicache/_3708_ ( .A(\myifu/myicache/_0103_ ), .Z(\myifu/myicache/_1705_ ) );
BUF_X1 \myifu/myicache/_3709_ ( .A(\myifu/myicache/_0104_ ), .Z(\myifu/myicache/_1706_ ) );
BUF_X1 \myifu/myicache/_3710_ ( .A(\myifu/myicache/_0105_ ), .Z(\myifu/myicache/_1707_ ) );
BUF_X1 \myifu/myicache/_3711_ ( .A(\myifu/myicache/_0106_ ), .Z(\myifu/myicache/_1708_ ) );
BUF_X1 \myifu/myicache/_3712_ ( .A(\myifu/myicache/_0107_ ), .Z(\myifu/myicache/_1709_ ) );
BUF_X1 \myifu/myicache/_3713_ ( .A(\myifu/myicache/_0108_ ), .Z(\myifu/myicache/_1710_ ) );
BUF_X1 \myifu/myicache/_3714_ ( .A(\myifu/myicache/_0109_ ), .Z(\myifu/myicache/_1711_ ) );
BUF_X1 \myifu/myicache/_3715_ ( .A(\myifu/myicache/_0110_ ), .Z(\myifu/myicache/_1712_ ) );
BUF_X1 \myifu/myicache/_3716_ ( .A(\myifu/myicache/_0111_ ), .Z(\myifu/myicache/_1713_ ) );
BUF_X1 \myifu/myicache/_3717_ ( .A(\myifu/myicache/_0112_ ), .Z(\myifu/myicache/_1714_ ) );
BUF_X1 \myifu/myicache/_3718_ ( .A(\myifu/myicache/_0113_ ), .Z(\myifu/myicache/_1715_ ) );
BUF_X1 \myifu/myicache/_3719_ ( .A(\myifu/myicache/_0114_ ), .Z(\myifu/myicache/_1716_ ) );
BUF_X1 \myifu/myicache/_3720_ ( .A(\myifu/myicache/_0115_ ), .Z(\myifu/myicache/_1717_ ) );
BUF_X1 \myifu/myicache/_3721_ ( .A(\myifu/myicache/_0116_ ), .Z(\myifu/myicache/_1718_ ) );
BUF_X1 \myifu/myicache/_3722_ ( .A(\myifu/myicache/_0117_ ), .Z(\myifu/myicache/_1719_ ) );
BUF_X1 \myifu/myicache/_3723_ ( .A(\myifu/myicache/_0118_ ), .Z(\myifu/myicache/_1720_ ) );
BUF_X1 \myifu/myicache/_3724_ ( .A(\myifu/myicache/_0119_ ), .Z(\myifu/myicache/_1721_ ) );
BUF_X1 \myifu/myicache/_3725_ ( .A(\myifu/myicache/_0120_ ), .Z(\myifu/myicache/_1722_ ) );
BUF_X1 \myifu/myicache/_3726_ ( .A(\myifu/myicache/_0121_ ), .Z(\myifu/myicache/_1723_ ) );
BUF_X1 \myifu/myicache/_3727_ ( .A(\myifu/myicache/_0122_ ), .Z(\myifu/myicache/_1724_ ) );
BUF_X1 \myifu/myicache/_3728_ ( .A(\myifu/myicache/_0123_ ), .Z(\myifu/myicache/_1725_ ) );
BUF_X1 \myifu/myicache/_3729_ ( .A(\myifu/myicache/_0124_ ), .Z(\myifu/myicache/_1726_ ) );
BUF_X1 \myifu/myicache/_3730_ ( .A(\myifu/myicache/_0125_ ), .Z(\myifu/myicache/_1727_ ) );
BUF_X1 \myifu/myicache/_3731_ ( .A(\myifu/myicache/_0126_ ), .Z(\myifu/myicache/_1728_ ) );
BUF_X1 \myifu/myicache/_3732_ ( .A(\myifu/myicache/_0127_ ), .Z(\myifu/myicache/_1729_ ) );
BUF_X1 \myifu/myicache/_3733_ ( .A(\myifu/myicache/_0128_ ), .Z(\myifu/myicache/_1730_ ) );
BUF_X1 \myifu/myicache/_3734_ ( .A(\myifu/myicache/_0129_ ), .Z(\myifu/myicache/_1731_ ) );
BUF_X1 \myifu/myicache/_3735_ ( .A(\myifu/myicache/_0130_ ), .Z(\myifu/myicache/_1732_ ) );
BUF_X1 \myifu/myicache/_3736_ ( .A(\myifu/myicache/_0131_ ), .Z(\myifu/myicache/_1733_ ) );
BUF_X1 \myifu/myicache/_3737_ ( .A(\myifu/myicache/_0132_ ), .Z(\myifu/myicache/_1734_ ) );
BUF_X1 \myifu/myicache/_3738_ ( .A(\myifu/myicache/_0133_ ), .Z(\myifu/myicache/_1735_ ) );
BUF_X1 \myifu/myicache/_3739_ ( .A(\myifu/myicache/_0134_ ), .Z(\myifu/myicache/_1736_ ) );
BUF_X1 \myifu/myicache/_3740_ ( .A(\myifu/myicache/_0135_ ), .Z(\myifu/myicache/_1737_ ) );
BUF_X1 \myifu/myicache/_3741_ ( .A(\myifu/myicache/_0136_ ), .Z(\myifu/myicache/_1738_ ) );
BUF_X1 \myifu/myicache/_3742_ ( .A(\myifu/myicache/_0137_ ), .Z(\myifu/myicache/_1739_ ) );
BUF_X1 \myifu/myicache/_3743_ ( .A(\myifu/myicache/_0138_ ), .Z(\myifu/myicache/_1740_ ) );
BUF_X1 \myifu/myicache/_3744_ ( .A(\myifu/myicache/_0139_ ), .Z(\myifu/myicache/_1741_ ) );
BUF_X1 \myifu/myicache/_3745_ ( .A(\myifu/myicache/_0140_ ), .Z(\myifu/myicache/_1742_ ) );
BUF_X1 \myifu/myicache/_3746_ ( .A(\myifu/myicache/_0141_ ), .Z(\myifu/myicache/_1743_ ) );
BUF_X1 \myifu/myicache/_3747_ ( .A(\myifu/myicache/_0142_ ), .Z(\myifu/myicache/_1744_ ) );
BUF_X1 \myifu/myicache/_3748_ ( .A(\myifu/myicache/_0143_ ), .Z(\myifu/myicache/_1745_ ) );
BUF_X1 \myifu/myicache/_3749_ ( .A(\myifu/myicache/_0144_ ), .Z(\myifu/myicache/_1746_ ) );
BUF_X1 \myifu/myicache/_3750_ ( .A(\myifu/myicache/_0145_ ), .Z(\myifu/myicache/_1747_ ) );
BUF_X1 \myifu/myicache/_3751_ ( .A(\myifu/myicache/_0146_ ), .Z(\myifu/myicache/_1748_ ) );
BUF_X1 \myifu/myicache/_3752_ ( .A(\myifu/myicache/_0147_ ), .Z(\myifu/myicache/_1749_ ) );
BUF_X1 \myifu/myicache/_3753_ ( .A(\myifu/myicache/_0148_ ), .Z(\myifu/myicache/_1750_ ) );
BUF_X1 \myifu/myicache/_3754_ ( .A(\myifu/myicache/_0149_ ), .Z(\myifu/myicache/_1751_ ) );
BUF_X1 \myifu/myicache/_3755_ ( .A(\myifu/myicache/_0150_ ), .Z(\myifu/myicache/_1752_ ) );
BUF_X1 \myifu/myicache/_3756_ ( .A(\myifu/myicache/_0151_ ), .Z(\myifu/myicache/_1753_ ) );
BUF_X1 \myifu/myicache/_3757_ ( .A(\myifu/myicache/_0152_ ), .Z(\myifu/myicache/_1754_ ) );
BUF_X1 \myifu/myicache/_3758_ ( .A(\myifu/myicache/_0153_ ), .Z(\myifu/myicache/_1755_ ) );
BUF_X1 \myifu/myicache/_3759_ ( .A(\myifu/myicache/_0154_ ), .Z(\myifu/myicache/_1756_ ) );
BUF_X1 \myifu/myicache/_3760_ ( .A(\myifu/myicache/_0155_ ), .Z(\myifu/myicache/_1757_ ) );
BUF_X1 \myifu/myicache/_3761_ ( .A(\myifu/myicache/_0156_ ), .Z(\myifu/myicache/_1758_ ) );
BUF_X1 \myifu/myicache/_3762_ ( .A(\myifu/myicache/_0157_ ), .Z(\myifu/myicache/_1759_ ) );
BUF_X1 \myifu/myicache/_3763_ ( .A(\myifu/myicache/_0158_ ), .Z(\myifu/myicache/_1760_ ) );
BUF_X1 \myifu/myicache/_3764_ ( .A(\myifu/myicache/_0159_ ), .Z(\myifu/myicache/_1761_ ) );
BUF_X1 \myifu/myicache/_3765_ ( .A(\myifu/myicache/_0160_ ), .Z(\myifu/myicache/_1762_ ) );
BUF_X1 \myifu/myicache/_3766_ ( .A(\myifu/myicache/_0161_ ), .Z(\myifu/myicache/_1763_ ) );
BUF_X1 \myifu/myicache/_3767_ ( .A(\myifu/myicache/_0162_ ), .Z(\myifu/myicache/_1764_ ) );
BUF_X1 \myifu/myicache/_3768_ ( .A(\myifu/myicache/_0163_ ), .Z(\myifu/myicache/_1765_ ) );
BUF_X1 \myifu/myicache/_3769_ ( .A(\myifu/myicache/_0164_ ), .Z(\myifu/myicache/_1766_ ) );
BUF_X1 \myifu/myicache/_3770_ ( .A(\myifu/myicache/_0165_ ), .Z(\myifu/myicache/_1767_ ) );
BUF_X1 \myifu/myicache/_3771_ ( .A(\myifu/myicache/_0166_ ), .Z(\myifu/myicache/_1768_ ) );
BUF_X1 \myifu/myicache/_3772_ ( .A(\myifu/myicache/_0167_ ), .Z(\myifu/myicache/_1769_ ) );
BUF_X1 \myifu/myicache/_3773_ ( .A(\myifu/myicache/_0168_ ), .Z(\myifu/myicache/_1770_ ) );
BUF_X1 \myifu/myicache/_3774_ ( .A(\myifu/myicache/_0169_ ), .Z(\myifu/myicache/_1771_ ) );
BUF_X1 \myifu/myicache/_3775_ ( .A(\myifu/myicache/_0170_ ), .Z(\myifu/myicache/_1772_ ) );
BUF_X1 \myifu/myicache/_3776_ ( .A(\myifu/myicache/_0171_ ), .Z(\myifu/myicache/_1773_ ) );
BUF_X1 \myifu/myicache/_3777_ ( .A(\myifu/myicache/_0172_ ), .Z(\myifu/myicache/_1774_ ) );
BUF_X1 \myifu/myicache/_3778_ ( .A(\myifu/myicache/_0173_ ), .Z(\myifu/myicache/_1775_ ) );
BUF_X1 \myifu/myicache/_3779_ ( .A(\myifu/myicache/_0174_ ), .Z(\myifu/myicache/_1776_ ) );
BUF_X1 \myifu/myicache/_3780_ ( .A(\myifu/myicache/_0175_ ), .Z(\myifu/myicache/_1777_ ) );
BUF_X1 \myifu/myicache/_3781_ ( .A(\myifu/myicache/_0176_ ), .Z(\myifu/myicache/_1778_ ) );
BUF_X1 \myifu/myicache/_3782_ ( .A(\myifu/myicache/_0177_ ), .Z(\myifu/myicache/_1779_ ) );
BUF_X1 \myifu/myicache/_3783_ ( .A(\myifu/myicache/_0178_ ), .Z(\myifu/myicache/_1780_ ) );
BUF_X1 \myifu/myicache/_3784_ ( .A(\myifu/myicache/_0179_ ), .Z(\myifu/myicache/_1781_ ) );
BUF_X1 \myifu/myicache/_3785_ ( .A(\myifu/myicache/_0180_ ), .Z(\myifu/myicache/_1782_ ) );
BUF_X1 \myifu/myicache/_3786_ ( .A(\myifu/myicache/_0181_ ), .Z(\myifu/myicache/_1783_ ) );
BUF_X1 \myifu/myicache/_3787_ ( .A(\myifu/myicache/_0182_ ), .Z(\myifu/myicache/_1784_ ) );
BUF_X1 \myifu/myicache/_3788_ ( .A(\myifu/myicache/_0183_ ), .Z(\myifu/myicache/_1785_ ) );
BUF_X1 \myifu/myicache/_3789_ ( .A(\myifu/myicache/_0184_ ), .Z(\myifu/myicache/_1786_ ) );
BUF_X1 \myifu/myicache/_3790_ ( .A(\myifu/myicache/_0185_ ), .Z(\myifu/myicache/_1787_ ) );
BUF_X1 \myifu/myicache/_3791_ ( .A(\myifu/myicache/_0186_ ), .Z(\myifu/myicache/_1788_ ) );
BUF_X1 \myifu/myicache/_3792_ ( .A(\myifu/myicache/_0187_ ), .Z(\myifu/myicache/_1789_ ) );
BUF_X1 \myifu/myicache/_3793_ ( .A(\myifu/myicache/_0188_ ), .Z(\myifu/myicache/_1790_ ) );
BUF_X1 \myifu/myicache/_3794_ ( .A(\myifu/myicache/_0189_ ), .Z(\myifu/myicache/_1791_ ) );
BUF_X1 \myifu/myicache/_3795_ ( .A(\myifu/myicache/_0190_ ), .Z(\myifu/myicache/_1792_ ) );
BUF_X1 \myifu/myicache/_3796_ ( .A(\myifu/myicache/_0191_ ), .Z(\myifu/myicache/_1793_ ) );
BUF_X1 \myifu/myicache/_3797_ ( .A(\myifu/myicache/_0192_ ), .Z(\myifu/myicache/_1794_ ) );
BUF_X1 \myifu/myicache/_3798_ ( .A(\myifu/myicache/_0193_ ), .Z(\myifu/myicache/_1795_ ) );
BUF_X1 \myifu/myicache/_3799_ ( .A(\myifu/myicache/_0194_ ), .Z(\myifu/myicache/_1796_ ) );
BUF_X1 \myifu/myicache/_3800_ ( .A(\myifu/myicache/_0195_ ), .Z(\myifu/myicache/_1797_ ) );
BUF_X1 \myifu/myicache/_3801_ ( .A(\myifu/myicache/_0196_ ), .Z(\myifu/myicache/_1798_ ) );
BUF_X1 \myifu/myicache/_3802_ ( .A(\myifu/myicache/_0197_ ), .Z(\myifu/myicache/_1799_ ) );
BUF_X1 \myifu/myicache/_3803_ ( .A(\myifu/myicache/_0198_ ), .Z(\myifu/myicache/_1800_ ) );
BUF_X1 \myifu/myicache/_3804_ ( .A(\myifu/myicache/_0199_ ), .Z(\myifu/myicache/_1801_ ) );
BUF_X1 \myifu/myicache/_3805_ ( .A(\myifu/myicache/_0200_ ), .Z(\myifu/myicache/_1802_ ) );
BUF_X1 \myifu/myicache/_3806_ ( .A(\myifu/myicache/_0201_ ), .Z(\myifu/myicache/_1803_ ) );
BUF_X1 \myifu/myicache/_3807_ ( .A(\myifu/myicache/_0202_ ), .Z(\myifu/myicache/_1804_ ) );
BUF_X1 \myifu/myicache/_3808_ ( .A(\myifu/myicache/_0203_ ), .Z(\myifu/myicache/_1805_ ) );
BUF_X1 \myifu/myicache/_3809_ ( .A(\myifu/myicache/_0204_ ), .Z(\myifu/myicache/_1806_ ) );
BUF_X1 \myifu/myicache/_3810_ ( .A(\myifu/myicache/_0205_ ), .Z(\myifu/myicache/_1807_ ) );
BUF_X1 \myifu/myicache/_3811_ ( .A(\myifu/myicache/_0206_ ), .Z(\myifu/myicache/_1808_ ) );
BUF_X1 \myifu/myicache/_3812_ ( .A(\myifu/myicache/_0207_ ), .Z(\myifu/myicache/_1809_ ) );
BUF_X1 \myifu/myicache/_3813_ ( .A(\myifu/myicache/_0208_ ), .Z(\myifu/myicache/_1810_ ) );
BUF_X1 \myifu/myicache/_3814_ ( .A(\myifu/myicache/_0209_ ), .Z(\myifu/myicache/_1811_ ) );
BUF_X1 \myifu/myicache/_3815_ ( .A(\myifu/myicache/_0210_ ), .Z(\myifu/myicache/_1812_ ) );
BUF_X1 \myifu/myicache/_3816_ ( .A(\myifu/myicache/_0211_ ), .Z(\myifu/myicache/_1813_ ) );
BUF_X1 \myifu/myicache/_3817_ ( .A(\myifu/myicache/_0212_ ), .Z(\myifu/myicache/_1814_ ) );
BUF_X1 \myifu/myicache/_3818_ ( .A(\myifu/myicache/_0213_ ), .Z(\myifu/myicache/_1815_ ) );
BUF_X1 \myifu/myicache/_3819_ ( .A(\myifu/myicache/_0214_ ), .Z(\myifu/myicache/_1816_ ) );
BUF_X1 \myifu/myicache/_3820_ ( .A(\myifu/myicache/_0215_ ), .Z(\myifu/myicache/_1817_ ) );
BUF_X1 \myifu/myicache/_3821_ ( .A(\myifu/myicache/_0216_ ), .Z(\myifu/myicache/_1818_ ) );
BUF_X1 \myifu/myicache/_3822_ ( .A(\myifu/myicache/_0217_ ), .Z(\myifu/myicache/_1819_ ) );
BUF_X1 \myifu/myicache/_3823_ ( .A(\myifu/myicache/_0218_ ), .Z(\myifu/myicache/_1820_ ) );
BUF_X1 \myifu/myicache/_3824_ ( .A(\myifu/myicache/_0219_ ), .Z(\myifu/myicache/_1821_ ) );
BUF_X1 \myifu/myicache/_3825_ ( .A(\myifu/myicache/_0220_ ), .Z(\myifu/myicache/_1822_ ) );
BUF_X1 \myifu/myicache/_3826_ ( .A(\myifu/myicache/_0221_ ), .Z(\myifu/myicache/_1823_ ) );
BUF_X1 \myifu/myicache/_3827_ ( .A(\myifu/myicache/_0222_ ), .Z(\myifu/myicache/_1824_ ) );
BUF_X1 \myifu/myicache/_3828_ ( .A(\myifu/myicache/_0223_ ), .Z(\myifu/myicache/_1825_ ) );
BUF_X1 \myifu/myicache/_3829_ ( .A(\myifu/myicache/_0224_ ), .Z(\myifu/myicache/_1826_ ) );
BUF_X1 \myifu/myicache/_3830_ ( .A(\myifu/myicache/_0225_ ), .Z(\myifu/myicache/_1827_ ) );
BUF_X1 \myifu/myicache/_3831_ ( .A(\myifu/myicache/_0226_ ), .Z(\myifu/myicache/_1828_ ) );
BUF_X1 \myifu/myicache/_3832_ ( .A(\araddr_IFU [5] ), .Z(\myifu/myicache/_1173_ ) );
BUF_X1 \myifu/myicache/_3833_ ( .A(\myifu/myicache/_0227_ ), .Z(\myifu/myicache/_1829_ ) );
BUF_X1 \myifu/myicache/_3834_ ( .A(\araddr_IFU [6] ), .Z(\myifu/myicache/_1184_ ) );
BUF_X1 \myifu/myicache/_3835_ ( .A(\myifu/myicache/_0228_ ), .Z(\myifu/myicache/_1830_ ) );
BUF_X1 \myifu/myicache/_3836_ ( .A(\araddr_IFU [7] ), .Z(\myifu/myicache/_1192_ ) );
BUF_X1 \myifu/myicache/_3837_ ( .A(\myifu/myicache/_0229_ ), .Z(\myifu/myicache/_1831_ ) );
BUF_X1 \myifu/myicache/_3838_ ( .A(\araddr_IFU [8] ), .Z(\myifu/myicache/_1193_ ) );
BUF_X1 \myifu/myicache/_3839_ ( .A(\myifu/myicache/_0230_ ), .Z(\myifu/myicache/_1832_ ) );
BUF_X1 \myifu/myicache/_3840_ ( .A(\araddr_IFU [9] ), .Z(\myifu/myicache/_1194_ ) );
BUF_X1 \myifu/myicache/_3841_ ( .A(\myifu/myicache/_0231_ ), .Z(\myifu/myicache/_1833_ ) );
BUF_X1 \myifu/myicache/_3842_ ( .A(\araddr_IFU [10] ), .Z(\myifu/myicache/_1195_ ) );
BUF_X1 \myifu/myicache/_3843_ ( .A(\myifu/myicache/_0232_ ), .Z(\myifu/myicache/_1834_ ) );
BUF_X1 \myifu/myicache/_3844_ ( .A(\araddr_IFU [11] ), .Z(\myifu/myicache/_1196_ ) );
BUF_X1 \myifu/myicache/_3845_ ( .A(\myifu/myicache/_0233_ ), .Z(\myifu/myicache/_1835_ ) );
BUF_X1 \myifu/myicache/_3846_ ( .A(\araddr_IFU [12] ), .Z(\myifu/myicache/_1197_ ) );
BUF_X1 \myifu/myicache/_3847_ ( .A(\myifu/myicache/_0234_ ), .Z(\myifu/myicache/_1836_ ) );
BUF_X1 \myifu/myicache/_3848_ ( .A(\araddr_IFU [13] ), .Z(\myifu/myicache/_1198_ ) );
BUF_X1 \myifu/myicache/_3849_ ( .A(\myifu/myicache/_0235_ ), .Z(\myifu/myicache/_1837_ ) );
BUF_X1 \myifu/myicache/_3850_ ( .A(\araddr_IFU [14] ), .Z(\myifu/myicache/_1199_ ) );
BUF_X1 \myifu/myicache/_3851_ ( .A(\myifu/myicache/_0236_ ), .Z(\myifu/myicache/_1838_ ) );
BUF_X1 \myifu/myicache/_3852_ ( .A(\araddr_IFU [15] ), .Z(\myifu/myicache/_1174_ ) );
BUF_X1 \myifu/myicache/_3853_ ( .A(\myifu/myicache/_0237_ ), .Z(\myifu/myicache/_1839_ ) );
BUF_X1 \myifu/myicache/_3854_ ( .A(\araddr_IFU [16] ), .Z(\myifu/myicache/_1175_ ) );
BUF_X1 \myifu/myicache/_3855_ ( .A(\myifu/myicache/_0238_ ), .Z(\myifu/myicache/_1840_ ) );
BUF_X1 \myifu/myicache/_3856_ ( .A(\araddr_IFU [17] ), .Z(\myifu/myicache/_1176_ ) );
BUF_X1 \myifu/myicache/_3857_ ( .A(\myifu/myicache/_0239_ ), .Z(\myifu/myicache/_1841_ ) );
BUF_X1 \myifu/myicache/_3858_ ( .A(\araddr_IFU [18] ), .Z(\myifu/myicache/_1177_ ) );
BUF_X1 \myifu/myicache/_3859_ ( .A(\myifu/myicache/_0240_ ), .Z(\myifu/myicache/_1842_ ) );
BUF_X1 \myifu/myicache/_3860_ ( .A(\araddr_IFU [19] ), .Z(\myifu/myicache/_1178_ ) );
BUF_X1 \myifu/myicache/_3861_ ( .A(\myifu/myicache/_0241_ ), .Z(\myifu/myicache/_1843_ ) );
BUF_X1 \myifu/myicache/_3862_ ( .A(\araddr_IFU [20] ), .Z(\myifu/myicache/_1179_ ) );
BUF_X1 \myifu/myicache/_3863_ ( .A(\myifu/myicache/_0242_ ), .Z(\myifu/myicache/_1844_ ) );
BUF_X1 \myifu/myicache/_3864_ ( .A(\araddr_IFU [21] ), .Z(\myifu/myicache/_1180_ ) );
BUF_X1 \myifu/myicache/_3865_ ( .A(\myifu/myicache/_0243_ ), .Z(\myifu/myicache/_1845_ ) );
BUF_X1 \myifu/myicache/_3866_ ( .A(\araddr_IFU [22] ), .Z(\myifu/myicache/_1181_ ) );
BUF_X1 \myifu/myicache/_3867_ ( .A(\myifu/myicache/_0244_ ), .Z(\myifu/myicache/_1846_ ) );
BUF_X1 \myifu/myicache/_3868_ ( .A(\araddr_IFU [23] ), .Z(\myifu/myicache/_1182_ ) );
BUF_X1 \myifu/myicache/_3869_ ( .A(\myifu/myicache/_0245_ ), .Z(\myifu/myicache/_1847_ ) );
BUF_X1 \myifu/myicache/_3870_ ( .A(\araddr_IFU [24] ), .Z(\myifu/myicache/_1183_ ) );
BUF_X1 \myifu/myicache/_3871_ ( .A(\myifu/myicache/_0246_ ), .Z(\myifu/myicache/_1848_ ) );
BUF_X1 \myifu/myicache/_3872_ ( .A(\araddr_IFU [25] ), .Z(\myifu/myicache/_1185_ ) );
BUF_X1 \myifu/myicache/_3873_ ( .A(\myifu/myicache/_0247_ ), .Z(\myifu/myicache/_1849_ ) );
BUF_X1 \myifu/myicache/_3874_ ( .A(\araddr_IFU [26] ), .Z(\myifu/myicache/_1186_ ) );
BUF_X1 \myifu/myicache/_3875_ ( .A(\myifu/myicache/_0248_ ), .Z(\myifu/myicache/_1850_ ) );
BUF_X1 \myifu/myicache/_3876_ ( .A(\araddr_IFU [27] ), .Z(\myifu/myicache/_1187_ ) );
BUF_X1 \myifu/myicache/_3877_ ( .A(\myifu/myicache/_0249_ ), .Z(\myifu/myicache/_1851_ ) );
BUF_X1 \myifu/myicache/_3878_ ( .A(\araddr_IFU [28] ), .Z(\myifu/myicache/_1188_ ) );
BUF_X1 \myifu/myicache/_3879_ ( .A(\myifu/myicache/_0250_ ), .Z(\myifu/myicache/_1852_ ) );
BUF_X1 \myifu/myicache/_3880_ ( .A(\araddr_IFU [29] ), .Z(\myifu/myicache/_1189_ ) );
BUF_X1 \myifu/myicache/_3881_ ( .A(\myifu/myicache/_0251_ ), .Z(\myifu/myicache/_1853_ ) );
BUF_X1 \myifu/myicache/_3882_ ( .A(\araddr_IFU [30] ), .Z(\myifu/myicache/_1190_ ) );
BUF_X1 \myifu/myicache/_3883_ ( .A(\myifu/myicache/_0252_ ), .Z(\myifu/myicache/_1854_ ) );
BUF_X1 \myifu/myicache/_3884_ ( .A(\araddr_IFU [31] ), .Z(\myifu/myicache/_1191_ ) );
BUF_X1 \myifu/myicache/_3885_ ( .A(\myifu/myicache/_0253_ ), .Z(\myifu/myicache/_1855_ ) );
BUF_X1 \myifu/myicache/_3886_ ( .A(\myifu/myicache/_0254_ ), .Z(\myifu/myicache/_1856_ ) );
BUF_X1 \myifu/myicache/_3887_ ( .A(\myifu/myicache/_0255_ ), .Z(\myifu/myicache/_1857_ ) );
BUF_X1 \myifu/myicache/_3888_ ( .A(\myifu/myicache/_0256_ ), .Z(\myifu/myicache/_1858_ ) );
BUF_X1 \myifu/myicache/_3889_ ( .A(\myifu/myicache/_0257_ ), .Z(\myifu/myicache/_1859_ ) );
BUF_X1 \myifu/myicache/_3890_ ( .A(\myifu/myicache/_0258_ ), .Z(\myifu/myicache/_1860_ ) );
BUF_X1 \myifu/myicache/_3891_ ( .A(\myifu/myicache/_0259_ ), .Z(\myifu/myicache/_1861_ ) );
BUF_X1 \myifu/myicache/_3892_ ( .A(\myifu/myicache/_0260_ ), .Z(\myifu/myicache/_1862_ ) );
BUF_X1 \myifu/myicache/_3893_ ( .A(\myifu/myicache/_0261_ ), .Z(\myifu/myicache/_1863_ ) );
BUF_X1 \myifu/myicache/_3894_ ( .A(\myifu/myicache/_0262_ ), .Z(\myifu/myicache/_1864_ ) );
BUF_X1 \myifu/myicache/_3895_ ( .A(\myifu/myicache/_0263_ ), .Z(\myifu/myicache/_1865_ ) );
BUF_X1 \myifu/myicache/_3896_ ( .A(\myifu/myicache/_0264_ ), .Z(\myifu/myicache/_1866_ ) );
BUF_X1 \myifu/myicache/_3897_ ( .A(\myifu/myicache/_0265_ ), .Z(\myifu/myicache/_1867_ ) );
BUF_X1 \myifu/myicache/_3898_ ( .A(\myifu/myicache/_0266_ ), .Z(\myifu/myicache/_1868_ ) );
BUF_X1 \myifu/myicache/_3899_ ( .A(\myifu/myicache/_0267_ ), .Z(\myifu/myicache/_1869_ ) );
BUF_X1 \myifu/myicache/_3900_ ( .A(\myifu/myicache/_0268_ ), .Z(\myifu/myicache/_1870_ ) );
BUF_X1 \myifu/myicache/_3901_ ( .A(\myifu/myicache/_0269_ ), .Z(\myifu/myicache/_1871_ ) );
BUF_X1 \myifu/myicache/_3902_ ( .A(\myifu/myicache/_0270_ ), .Z(\myifu/myicache/_1872_ ) );
BUF_X1 \myifu/myicache/_3903_ ( .A(\myifu/myicache/_0271_ ), .Z(\myifu/myicache/_1873_ ) );
BUF_X1 \myifu/myicache/_3904_ ( .A(\myifu/myicache/_0272_ ), .Z(\myifu/myicache/_1874_ ) );
BUF_X1 \myifu/myicache/_3905_ ( .A(\myifu/myicache/_0273_ ), .Z(\myifu/myicache/_1875_ ) );
BUF_X1 \myifu/myicache/_3906_ ( .A(\myifu/myicache/_0274_ ), .Z(\myifu/myicache/_1876_ ) );
BUF_X1 \myifu/myicache/_3907_ ( .A(\myifu/myicache/_0275_ ), .Z(\myifu/myicache/_1877_ ) );
BUF_X1 \myifu/myicache/_3908_ ( .A(\myifu/myicache/_0276_ ), .Z(\myifu/myicache/_1878_ ) );
BUF_X1 \myifu/myicache/_3909_ ( .A(\myifu/myicache/_0277_ ), .Z(\myifu/myicache/_1879_ ) );
BUF_X1 \myifu/myicache/_3910_ ( .A(\myifu/myicache/_0278_ ), .Z(\myifu/myicache/_1880_ ) );
BUF_X1 \myifu/myicache/_3911_ ( .A(\myifu/myicache/_0279_ ), .Z(\myifu/myicache/_1881_ ) );
BUF_X1 \myifu/myicache/_3912_ ( .A(\myifu/myicache/_0280_ ), .Z(\myifu/myicache/_1882_ ) );
BUF_X1 \myifu/myicache/_3913_ ( .A(\myifu/myicache/_0281_ ), .Z(\myifu/myicache/_1883_ ) );
BUF_X1 \myifu/myicache/_3914_ ( .A(\myifu/myicache/_0282_ ), .Z(\myifu/myicache/_1884_ ) );
BUF_X1 \myifu/myicache/_3915_ ( .A(\myifu/myicache/_0283_ ), .Z(\myifu/myicache/_1885_ ) );
BUF_X1 \myifu/myicache/_3916_ ( .A(\myifu/myicache/_0284_ ), .Z(\myifu/myicache/_1886_ ) );
BUF_X1 \myifu/myicache/_3917_ ( .A(\myifu/myicache/_0285_ ), .Z(\myifu/myicache/_1887_ ) );
BUF_X1 \myifu/myicache/_3918_ ( .A(\myifu/myicache/_0286_ ), .Z(\myifu/myicache/_1888_ ) );
BUF_X1 \myifu/myicache/_3919_ ( .A(\myifu/myicache/_0287_ ), .Z(\myifu/myicache/_1889_ ) );
BUF_X1 \myifu/myicache/_3920_ ( .A(\myifu/myicache/_0288_ ), .Z(\myifu/myicache/_1890_ ) );
BUF_X1 \myifu/myicache/_3921_ ( .A(\myifu/myicache/_0289_ ), .Z(\myifu/myicache/_1891_ ) );
BUF_X1 \myifu/myicache/_3922_ ( .A(\myifu/myicache/_0290_ ), .Z(\myifu/myicache/_1892_ ) );
BUF_X1 \myifu/myicache/_3923_ ( .A(\myifu/myicache/_0291_ ), .Z(\myifu/myicache/_1893_ ) );
BUF_X1 \myifu/myicache/_3924_ ( .A(\myifu/myicache/_0292_ ), .Z(\myifu/myicache/_1894_ ) );
BUF_X1 \myifu/myicache/_3925_ ( .A(\myifu/myicache/_0293_ ), .Z(\myifu/myicache/_1895_ ) );
BUF_X1 \myifu/myicache/_3926_ ( .A(\myifu/myicache/_0294_ ), .Z(\myifu/myicache/_1896_ ) );
BUF_X1 \myifu/myicache/_3927_ ( .A(\myifu/myicache/_0295_ ), .Z(\myifu/myicache/_1897_ ) );
BUF_X1 \myifu/myicache/_3928_ ( .A(\myifu/myicache/_0296_ ), .Z(\myifu/myicache/_1898_ ) );
BUF_X1 \myifu/myicache/_3929_ ( .A(\myifu/myicache/_0297_ ), .Z(\myifu/myicache/_1899_ ) );
BUF_X1 \myifu/myicache/_3930_ ( .A(\myifu/myicache/_0298_ ), .Z(\myifu/myicache/_1900_ ) );
BUF_X1 \myifu/myicache/_3931_ ( .A(\myifu/myicache/_0299_ ), .Z(\myifu/myicache/_1901_ ) );
BUF_X1 \myifu/myicache/_3932_ ( .A(\myifu/myicache/_0300_ ), .Z(\myifu/myicache/_1902_ ) );
BUF_X1 \myifu/myicache/_3933_ ( .A(\myifu/myicache/_0301_ ), .Z(\myifu/myicache/_1903_ ) );
BUF_X1 \myifu/myicache/_3934_ ( .A(\myifu/myicache/_0302_ ), .Z(\myifu/myicache/_1904_ ) );
BUF_X1 \myifu/myicache/_3935_ ( .A(\myifu/myicache/_0303_ ), .Z(\myifu/myicache/_1905_ ) );
BUF_X1 \myifu/myicache/_3936_ ( .A(\myifu/myicache/_0304_ ), .Z(\myifu/myicache/_1906_ ) );
BUF_X1 \myifu/myicache/_3937_ ( .A(\myifu/myicache/_0305_ ), .Z(\myifu/myicache/_1907_ ) );
BUF_X1 \myifu/myicache/_3938_ ( .A(\myifu/myicache/_0306_ ), .Z(\myifu/myicache/_1908_ ) );
BUF_X1 \myifu/myicache/_3939_ ( .A(\myifu/myicache/_0307_ ), .Z(\myifu/myicache/_1909_ ) );
BUF_X1 \myifu/myicache/_3940_ ( .A(\myifu/myicache/_0308_ ), .Z(\myifu/myicache/_1910_ ) );
BUF_X1 \myifu/myicache/_3941_ ( .A(\myifu/myicache/_0309_ ), .Z(\myifu/myicache/_1911_ ) );
BUF_X1 \myifu/myicache/_3942_ ( .A(\myifu/myicache/_0310_ ), .Z(\myifu/myicache/_1912_ ) );
BUF_X1 \myifu/myicache/_3943_ ( .A(\myifu/myicache/_0311_ ), .Z(\myifu/myicache/_1913_ ) );
BUF_X1 \myifu/myicache/_3944_ ( .A(\myifu/myicache/_0312_ ), .Z(\myifu/myicache/_1914_ ) );
BUF_X1 \myifu/myicache/_3945_ ( .A(\myifu/myicache/_0313_ ), .Z(\myifu/myicache/_1915_ ) );
BUF_X1 \myifu/myicache/_3946_ ( .A(\myifu/myicache/_0314_ ), .Z(\myifu/myicache/_1916_ ) );
BUF_X1 \myifu/myicache/_3947_ ( .A(\myifu/myicache/_0315_ ), .Z(\myifu/myicache/_1917_ ) );
BUF_X1 \myifu/myicache/_3948_ ( .A(\myifu/myicache/_0316_ ), .Z(\myifu/myicache/_1918_ ) );
BUF_X1 \myifu/myicache/_3949_ ( .A(\myifu/myicache/_0317_ ), .Z(\myifu/myicache/_1919_ ) );
BUF_X1 \myifu/myicache/_3950_ ( .A(\myifu/myicache/_0318_ ), .Z(\myifu/myicache/_1920_ ) );
BUF_X1 \myifu/myicache/_3951_ ( .A(\myifu/myicache/_0319_ ), .Z(\myifu/myicache/_1921_ ) );
BUF_X1 \myifu/myicache/_3952_ ( .A(\myifu/myicache/_0320_ ), .Z(\myifu/myicache/_1922_ ) );
BUF_X1 \myifu/myicache/_3953_ ( .A(\myifu/myicache/_0321_ ), .Z(\myifu/myicache/_1923_ ) );
BUF_X1 \myifu/myicache/_3954_ ( .A(\myifu/myicache/_0322_ ), .Z(\myifu/myicache/_1924_ ) );
BUF_X1 \myifu/myicache/_3955_ ( .A(\myifu/myicache/_0323_ ), .Z(\myifu/myicache/_1925_ ) );
BUF_X1 \myifu/myicache/_3956_ ( .A(\myifu/myicache/_0324_ ), .Z(\myifu/myicache/_1926_ ) );
BUF_X1 \myifu/myicache/_3957_ ( .A(\myifu/myicache/_0325_ ), .Z(\myifu/myicache/_1927_ ) );
BUF_X1 \myifu/myicache/_3958_ ( .A(\myifu/myicache/_0326_ ), .Z(\myifu/myicache/_1928_ ) );
BUF_X1 \myifu/myicache/_3959_ ( .A(\myifu/myicache/_0327_ ), .Z(\myifu/myicache/_1929_ ) );
BUF_X1 \myifu/myicache/_3960_ ( .A(\myifu/myicache/_0328_ ), .Z(\myifu/myicache/_1930_ ) );
BUF_X1 \myifu/myicache/_3961_ ( .A(\myifu/myicache/_0329_ ), .Z(\myifu/myicache/_1931_ ) );
BUF_X1 \myifu/myicache/_3962_ ( .A(\myifu/myicache/_0330_ ), .Z(\myifu/myicache/_1932_ ) );
BUF_X1 \myifu/myicache/_3963_ ( .A(\myifu/myicache/_0331_ ), .Z(\myifu/myicache/_1933_ ) );
BUF_X1 \myifu/myicache/_3964_ ( .A(\myifu/myicache/_0332_ ), .Z(\myifu/myicache/_1934_ ) );
BUF_X1 \myifu/myicache/_3965_ ( .A(\myifu/myicache/_0333_ ), .Z(\myifu/myicache/_1935_ ) );
BUF_X1 \myifu/myicache/_3966_ ( .A(\myifu/myicache/_0334_ ), .Z(\myifu/myicache/_1936_ ) );
BUF_X1 \myifu/myicache/_3967_ ( .A(\myifu/myicache/_0335_ ), .Z(\myifu/myicache/_1937_ ) );
BUF_X1 \myifu/myicache/_3968_ ( .A(\myifu/myicache/_0336_ ), .Z(\myifu/myicache/_1938_ ) );
BUF_X1 \myifu/myicache/_3969_ ( .A(\myifu/myicache/_0337_ ), .Z(\myifu/myicache/_1939_ ) );
BUF_X1 \myifu/myicache/_3970_ ( .A(\myifu/myicache/_0338_ ), .Z(\myifu/myicache/_1940_ ) );
BUF_X1 \myifu/myicache/_3971_ ( .A(\myifu/myicache/_0339_ ), .Z(\myifu/myicache/_1941_ ) );
BUF_X1 \myifu/myicache/_3972_ ( .A(\myifu/myicache/_0340_ ), .Z(\myifu/myicache/_1942_ ) );
BUF_X1 \myifu/myicache/_3973_ ( .A(\myifu/myicache/_0341_ ), .Z(\myifu/myicache/_1943_ ) );
BUF_X1 \myifu/myicache/_3974_ ( .A(\myifu/myicache/_0342_ ), .Z(\myifu/myicache/_1944_ ) );
BUF_X1 \myifu/myicache/_3975_ ( .A(\myifu/myicache/_0343_ ), .Z(\myifu/myicache/_1945_ ) );
BUF_X1 \myifu/myicache/_3976_ ( .A(\myifu/myicache/_0344_ ), .Z(\myifu/myicache/_1946_ ) );
BUF_X1 \myifu/myicache/_3977_ ( .A(\myifu/myicache/_0345_ ), .Z(\myifu/myicache/_1947_ ) );
BUF_X1 \myifu/myicache/_3978_ ( .A(\myifu/myicache/_0346_ ), .Z(\myifu/myicache/_1948_ ) );
BUF_X1 \myifu/myicache/_3979_ ( .A(\myifu/myicache/_0347_ ), .Z(\myifu/myicache/_1949_ ) );
BUF_X1 \myifu/myicache/_3980_ ( .A(\myifu/myicache/_0348_ ), .Z(\myifu/myicache/_1950_ ) );
BUF_X1 \myifu/myicache/_3981_ ( .A(\myifu/myicache/_0349_ ), .Z(\myifu/myicache/_1951_ ) );
BUF_X1 \myifu/myicache/_3982_ ( .A(\myifu/myicache/_0350_ ), .Z(\myifu/myicache/_1952_ ) );
BUF_X1 \myifu/myicache/_3983_ ( .A(\myifu/myicache/_0351_ ), .Z(\myifu/myicache/_1953_ ) );
BUF_X1 \myifu/myicache/_3984_ ( .A(\myifu/myicache/_0352_ ), .Z(\myifu/myicache/_1954_ ) );
BUF_X1 \myifu/myicache/_3985_ ( .A(\myifu/myicache/_0353_ ), .Z(\myifu/myicache/_1955_ ) );
BUF_X1 \myifu/myicache/_3986_ ( .A(\myifu/myicache/_0354_ ), .Z(\myifu/myicache/_1956_ ) );
BUF_X1 \myifu/myicache/_3987_ ( .A(\myifu/myicache/_0355_ ), .Z(\myifu/myicache/_1957_ ) );
BUF_X1 \myifu/myicache/_3988_ ( .A(\myifu/myicache/_0356_ ), .Z(\myifu/myicache/_1958_ ) );
BUF_X1 \myifu/myicache/_3989_ ( .A(\myifu/myicache/_0357_ ), .Z(\myifu/myicache/_1959_ ) );
BUF_X1 \myifu/myicache/_3990_ ( .A(\myifu/myicache/_0358_ ), .Z(\myifu/myicache/_1960_ ) );
BUF_X1 \myifu/myicache/_3991_ ( .A(\myifu/myicache/_0359_ ), .Z(\myifu/myicache/_1961_ ) );
BUF_X1 \myifu/myicache/_3992_ ( .A(\myifu/myicache/_0360_ ), .Z(\myifu/myicache/_1962_ ) );
BUF_X1 \myifu/myicache/_3993_ ( .A(\myifu/myicache/_0361_ ), .Z(\myifu/myicache/_1963_ ) );
BUF_X1 \myifu/myicache/_3994_ ( .A(\myifu/myicache/_0362_ ), .Z(\myifu/myicache/_1964_ ) );
BUF_X1 \myifu/myicache/_3995_ ( .A(\myifu/myicache/_0363_ ), .Z(\myifu/myicache/_1965_ ) );
BUF_X1 \myifu/myicache/_3996_ ( .A(\myifu/myicache/_0364_ ), .Z(\myifu/myicache/_1966_ ) );
BUF_X1 \myifu/myicache/_3997_ ( .A(\myifu/myicache/_0365_ ), .Z(\myifu/myicache/_1967_ ) );
BUF_X1 \myifu/myicache/_3998_ ( .A(\myifu/myicache/_0366_ ), .Z(\myifu/myicache/_1968_ ) );
BUF_X1 \myifu/myicache/_3999_ ( .A(\myifu/myicache/_0367_ ), .Z(\myifu/myicache/_1969_ ) );
INV_X2 \mylsu/_1366_ ( .A(fanout_net_26 ), .ZN(\mylsu/_0531_ ) );
INV_X1 \mylsu/_1367_ ( .A(\mylsu/_0298_ ), .ZN(\mylsu/_0532_ ) );
NAND3_X1 \mylsu/_1368_ ( .A1(\mylsu/_0531_ ), .A2(\mylsu/_0532_ ), .A3(\mylsu/_0917_ ), .ZN(\mylsu/_0533_ ) );
INV_X1 \mylsu/_1369_ ( .A(\mylsu/_0924_ ), .ZN(\mylsu/_0534_ ) );
NOR2_X1 \mylsu/_1370_ ( .A1(\mylsu/_0534_ ), .A2(\mylsu/_0925_ ), .ZN(\mylsu/_0535_ ) );
INV_X1 \mylsu/_1371_ ( .A(\mylsu/_0923_ ), .ZN(\mylsu/_0536_ ) );
AND2_X1 \mylsu/_1372_ ( .A1(\mylsu/_0535_ ), .A2(\mylsu/_0536_ ), .ZN(\mylsu/_0537_ ) );
AND4_X1 \mylsu/_1373_ ( .A1(\mylsu/_0929_ ), .A2(\mylsu/_0531_ ), .A3(\mylsu/_0532_ ), .A4(\mylsu/_1047_ ), .ZN(\mylsu/_0538_ ) );
INV_X1 \mylsu/_1374_ ( .A(\mylsu/_1047_ ), .ZN(\mylsu/_0539_ ) );
OAI211_X2 \mylsu/_1375_ ( .A(\mylsu/_0537_ ), .B(\mylsu/_0538_ ), .C1(\mylsu/_0539_ ), .C2(\mylsu/_0532_ ), .ZN(\mylsu/_0540_ ) );
INV_X1 \mylsu/_1376_ ( .A(\mylsu/_0913_ ), .ZN(\mylsu/_0541_ ) );
OAI21_X1 \mylsu/_1377_ ( .A(\mylsu/_0533_ ), .B1(\mylsu/_0540_ ), .B2(\mylsu/_0541_ ), .ZN(\mylsu/_0011_ ) );
INV_X1 \mylsu/_1378_ ( .A(\mylsu/_0904_ ), .ZN(\mylsu/_0542_ ) );
NOR4_X2 \mylsu/_1379_ ( .A1(\mylsu/_0542_ ), .A2(\mylsu/_0903_ ), .A3(\mylsu/_0906_ ), .A4(\mylsu/_0905_ ), .ZN(\mylsu/_0543_ ) );
NAND2_X1 \mylsu/_1380_ ( .A1(\mylsu/_0912_ ), .A2(\mylsu/_0907_ ), .ZN(\mylsu/_0544_ ) );
NOR3_X1 \mylsu/_1381_ ( .A1(\mylsu/_0544_ ), .A2(\mylsu/_0910_ ), .A3(\mylsu/_0909_ ), .ZN(\mylsu/_0545_ ) );
AND2_X4 \mylsu/_1382_ ( .A1(\mylsu/_0543_ ), .A2(\mylsu/_0545_ ), .ZN(\mylsu/_0546_ ) );
INV_X1 \mylsu/_1383_ ( .A(fanout_net_27 ), .ZN(\mylsu/_0547_ ) );
OR2_X4 \mylsu/_1384_ ( .A1(\mylsu/_0546_ ), .A2(\mylsu/_0547_ ), .ZN(\mylsu/_0548_ ) );
AND2_X4 \mylsu/_1385_ ( .A1(\mylsu/_0913_ ), .A2(\mylsu/_0929_ ), .ZN(\mylsu/_0549_ ) );
AND2_X1 \mylsu/_1386_ ( .A1(\mylsu/_0923_ ), .A2(\mylsu/_0924_ ), .ZN(\mylsu/_0550_ ) );
INV_X1 \mylsu/_1387_ ( .A(\mylsu/_0925_ ), .ZN(\mylsu/_0551_ ) );
NAND4_X1 \mylsu/_1388_ ( .A1(\mylsu/_0549_ ), .A2(\mylsu/_0550_ ), .A3(\mylsu/_0551_ ), .A4(\mylsu/_0078_ ), .ZN(\mylsu/_0552_ ) );
AOI21_X1 \mylsu/_1389_ ( .A(fanout_net_26 ), .B1(\mylsu/_0548_ ), .B2(\mylsu/_0552_ ), .ZN(\mylsu/_0010_ ) );
INV_X1 \mylsu/_1390_ ( .A(\mylsu/_0303_ ), .ZN(\mylsu/_0553_ ) );
OR3_X1 \mylsu/_1391_ ( .A1(\mylsu/_0553_ ), .A2(\mylsu/_0308_ ), .A3(\mylsu/_0305_ ), .ZN(\mylsu/_0554_ ) );
INV_X1 \mylsu/_1392_ ( .A(\mylsu/_0307_ ), .ZN(\mylsu/_0555_ ) );
INV_X1 \mylsu/_1393_ ( .A(\mylsu/_0304_ ), .ZN(\mylsu/_0556_ ) );
NAND4_X1 \mylsu/_1394_ ( .A1(\mylsu/_0555_ ), .A2(\mylsu/_0556_ ), .A3(\mylsu/_0309_ ), .A4(\mylsu/_0302_ ), .ZN(\mylsu/_0557_ ) );
NOR2_X1 \mylsu/_1395_ ( .A1(\mylsu/_0554_ ), .A2(\mylsu/_0557_ ), .ZN(\mylsu/_0558_ ) );
AOI22_X1 \mylsu/_1396_ ( .A1(\mylsu/_0546_ ), .A2(fanout_net_27 ), .B1(\mylsu/_0558_ ), .B2(\mylsu/_0914_ ), .ZN(\mylsu/_0559_ ) );
OAI211_X2 \mylsu/_1397_ ( .A(\mylsu/_0535_ ), .B(\mylsu/_0929_ ), .C1(\mylsu/_0536_ ), .C2(\mylsu/_0078_ ), .ZN(\mylsu/_0560_ ) );
NOR2_X1 \mylsu/_1398_ ( .A1(\mylsu/_1047_ ), .A2(\mylsu/_0298_ ), .ZN(\mylsu/_0561_ ) );
AOI21_X1 \mylsu/_1399_ ( .A(\mylsu/_0560_ ), .B1(\mylsu/_0537_ ), .B2(\mylsu/_0561_ ), .ZN(\mylsu/_0562_ ) );
OAI211_X2 \mylsu/_1400_ ( .A(\mylsu/_0559_ ), .B(\mylsu/_0531_ ), .C1(\mylsu/_0541_ ), .C2(\mylsu/_0562_ ), .ZN(\mylsu/_0007_ ) );
INV_X1 \mylsu/_1401_ ( .A(\mylsu/_0914_ ), .ZN(\mylsu/_0563_ ) );
NOR2_X1 \mylsu/_1402_ ( .A1(\mylsu/_0558_ ), .A2(\mylsu/_0563_ ), .ZN(\mylsu/_0564_ ) );
AOI21_X1 \mylsu/_1403_ ( .A(\mylsu/_0564_ ), .B1(\mylsu/_0298_ ), .B2(\mylsu/_0917_ ), .ZN(\mylsu/_0565_ ) );
AND2_X1 \mylsu/_1404_ ( .A1(\mylsu/_0549_ ), .A2(\mylsu/_0531_ ), .ZN(\mylsu/_0566_ ) );
BUF_X4 \mylsu/_1405_ ( .A(\mylsu/_0566_ ), .Z(\mylsu/_0567_ ) );
AND3_X1 \mylsu/_1406_ ( .A1(\mylsu/_0537_ ), .A2(\mylsu/_0298_ ), .A3(\mylsu/_0567_ ), .ZN(\mylsu/_0568_ ) );
AOI21_X1 \mylsu/_1407_ ( .A(\mylsu/_0568_ ), .B1(\mylsu/_0531_ ), .B2(\mylsu/_0915_ ), .ZN(\mylsu/_0569_ ) );
OAI22_X1 \mylsu/_1408_ ( .A1(fanout_net_26 ), .A2(\mylsu/_0565_ ), .B1(\mylsu/_0569_ ), .B2(\mylsu/_0539_ ), .ZN(\mylsu/_0008_ ) );
INV_X1 \mylsu/_1409_ ( .A(\mylsu/_0568_ ), .ZN(\mylsu/_0570_ ) );
NAND3_X1 \mylsu/_1410_ ( .A1(\mylsu/_0531_ ), .A2(\mylsu/_0539_ ), .A3(\mylsu/_0915_ ), .ZN(\mylsu/_0571_ ) );
AOI22_X1 \mylsu/_1411_ ( .A1(\mylsu/_0570_ ), .A2(\mylsu/_0571_ ), .B1(\mylsu/_1047_ ), .B2(\mylsu/_0298_ ), .ZN(\mylsu/_0009_ ) );
OR4_X1 \mylsu/_1412_ ( .A1(\mylsu/_0536_ ), .A2(\mylsu/_0534_ ), .A3(\mylsu/_0925_ ), .A4(\mylsu/_0012_ ), .ZN(\mylsu/_0572_ ) );
INV_X1 \mylsu/_1413_ ( .A(\mylsu/_0929_ ), .ZN(\mylsu/_0573_ ) );
NOR2_X2 \mylsu/_1414_ ( .A1(\mylsu/_0572_ ), .A2(\mylsu/_0573_ ), .ZN(\mylsu/_0574_ ) );
BUF_X4 \mylsu/_1415_ ( .A(\mylsu/_0574_ ), .Z(\mylsu/_0079_ ) );
BUF_X2 \mylsu/_1416_ ( .A(\mylsu/_0547_ ), .Z(\mylsu/_0575_ ) );
OAI21_X1 \mylsu/_1417_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0572_ ), .B2(\mylsu/_0573_ ), .ZN(\mylsu/_0908_ ) );
NOR4_X1 \mylsu/_1418_ ( .A1(\mylsu/_0534_ ), .A2(\mylsu/_0923_ ), .A3(\mylsu/_0925_ ), .A4(\mylsu/_0012_ ), .ZN(\mylsu/_0576_ ) );
NAND2_X2 \mylsu/_1419_ ( .A1(\mylsu/_0576_ ), .A2(\mylsu/_0929_ ), .ZN(\mylsu/_0577_ ) );
BUF_X4 \mylsu/_1420_ ( .A(\mylsu/_0577_ ), .Z(\mylsu/_0578_ ) );
INV_X1 \mylsu/_1421_ ( .A(\mylsu/_0917_ ), .ZN(\mylsu/_0579_ ) );
NAND2_X1 \mylsu/_1422_ ( .A1(\mylsu/_0578_ ), .A2(\mylsu/_0579_ ), .ZN(\mylsu/_0301_ ) );
INV_X1 \mylsu/_1423_ ( .A(\mylsu/_0915_ ), .ZN(\mylsu/_0580_ ) );
NAND2_X1 \mylsu/_1424_ ( .A1(\mylsu/_0578_ ), .A2(\mylsu/_0580_ ), .ZN(\mylsu/_1052_ ) );
NAND4_X1 \mylsu/_1425_ ( .A1(\mylsu/_0578_ ), .A2(\mylsu/_0563_ ), .A3(\mylsu/_0579_ ), .A4(\mylsu/_0580_ ), .ZN(\mylsu/_0306_ ) );
NAND2_X1 \mylsu/_1426_ ( .A1(\mylsu/_0541_ ), .A2(\mylsu/_0579_ ), .ZN(\mylsu/_0838_ ) );
MUX2_X1 \mylsu/_1427_ ( .A(\mylsu/_0046_ ), .B(fanout_net_25 ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0014_ ) );
MUX2_X1 \mylsu/_1428_ ( .A(\mylsu/_0057_ ), .B(\mylsu/_0321_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0025_ ) );
MUX2_X1 \mylsu/_1429_ ( .A(\mylsu/_0068_ ), .B(\mylsu/_0332_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0036_ ) );
MUX2_X1 \mylsu/_1430_ ( .A(\mylsu/_0071_ ), .B(\mylsu/_0335_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0039_ ) );
MUX2_X1 \mylsu/_1431_ ( .A(\mylsu/_0072_ ), .B(\mylsu/_0336_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0040_ ) );
MUX2_X1 \mylsu/_1432_ ( .A(\mylsu/_0073_ ), .B(\mylsu/_0337_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0041_ ) );
MUX2_X1 \mylsu/_1433_ ( .A(\mylsu/_0074_ ), .B(\mylsu/_0338_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0042_ ) );
MUX2_X1 \mylsu/_1434_ ( .A(\mylsu/_0075_ ), .B(\mylsu/_0339_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0043_ ) );
MUX2_X1 \mylsu/_1435_ ( .A(\mylsu/_0076_ ), .B(\mylsu/_0340_ ), .S(\mylsu/_0079_ ), .Z(\mylsu/_0044_ ) );
BUF_X4 \mylsu/_1436_ ( .A(\mylsu/_0574_ ), .Z(\mylsu/_0581_ ) );
MUX2_X1 \mylsu/_1437_ ( .A(\mylsu/_0077_ ), .B(\mylsu/_0341_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0045_ ) );
MUX2_X1 \mylsu/_1438_ ( .A(\mylsu/_0047_ ), .B(\mylsu/_0311_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0015_ ) );
MUX2_X1 \mylsu/_1439_ ( .A(\mylsu/_0048_ ), .B(\mylsu/_0312_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0016_ ) );
MUX2_X1 \mylsu/_1440_ ( .A(\mylsu/_0049_ ), .B(\mylsu/_0313_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0017_ ) );
MUX2_X1 \mylsu/_1441_ ( .A(\mylsu/_0050_ ), .B(\mylsu/_0314_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0018_ ) );
MUX2_X1 \mylsu/_1442_ ( .A(\mylsu/_0051_ ), .B(\mylsu/_0315_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0019_ ) );
MUX2_X1 \mylsu/_1443_ ( .A(\mylsu/_0052_ ), .B(\mylsu/_0316_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0020_ ) );
MUX2_X1 \mylsu/_1444_ ( .A(\mylsu/_0053_ ), .B(\mylsu/_0317_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0021_ ) );
MUX2_X1 \mylsu/_1445_ ( .A(\mylsu/_0054_ ), .B(\mylsu/_0318_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0022_ ) );
MUX2_X1 \mylsu/_1446_ ( .A(\mylsu/_0055_ ), .B(\mylsu/_0319_ ), .S(\mylsu/_0581_ ), .Z(\mylsu/_0023_ ) );
BUF_X4 \mylsu/_1447_ ( .A(\mylsu/_0574_ ), .Z(\mylsu/_0582_ ) );
MUX2_X1 \mylsu/_1448_ ( .A(\mylsu/_0056_ ), .B(\mylsu/_0320_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0024_ ) );
MUX2_X1 \mylsu/_1449_ ( .A(\mylsu/_0058_ ), .B(\mylsu/_0322_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0026_ ) );
MUX2_X1 \mylsu/_1450_ ( .A(\mylsu/_0059_ ), .B(\mylsu/_0323_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0027_ ) );
MUX2_X1 \mylsu/_1451_ ( .A(\mylsu/_0060_ ), .B(\mylsu/_0324_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0028_ ) );
MUX2_X1 \mylsu/_1452_ ( .A(\mylsu/_0061_ ), .B(\mylsu/_0325_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0029_ ) );
MUX2_X1 \mylsu/_1453_ ( .A(\mylsu/_0062_ ), .B(\mylsu/_0326_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0030_ ) );
MUX2_X1 \mylsu/_1454_ ( .A(\mylsu/_0063_ ), .B(\mylsu/_0327_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0031_ ) );
MUX2_X1 \mylsu/_1455_ ( .A(\mylsu/_0064_ ), .B(\mylsu/_0328_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0032_ ) );
MUX2_X1 \mylsu/_1456_ ( .A(\mylsu/_0065_ ), .B(\mylsu/_0329_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0033_ ) );
MUX2_X1 \mylsu/_1457_ ( .A(\mylsu/_0066_ ), .B(\mylsu/_0330_ ), .S(\mylsu/_0582_ ), .Z(\mylsu/_0034_ ) );
MUX2_X1 \mylsu/_1458_ ( .A(\mylsu/_0067_ ), .B(\mylsu/_0331_ ), .S(\mylsu/_0574_ ), .Z(\mylsu/_0035_ ) );
MUX2_X1 \mylsu/_1459_ ( .A(\mylsu/_0069_ ), .B(\mylsu/_0333_ ), .S(\mylsu/_0574_ ), .Z(\mylsu/_0037_ ) );
MUX2_X1 \mylsu/_1460_ ( .A(\mylsu/_0070_ ), .B(\mylsu/_0334_ ), .S(\mylsu/_0574_ ), .Z(\mylsu/_0038_ ) );
INV_X1 \mylsu/_1461_ ( .A(\mylsu/_0918_ ), .ZN(\mylsu/_0583_ ) );
NOR4_X1 \mylsu/_1462_ ( .A1(\mylsu/_0583_ ), .A2(\mylsu/_0921_ ), .A3(\mylsu/_0920_ ), .A4(\mylsu/_0922_ ), .ZN(\mylsu/_0584_ ) );
AND4_X1 \mylsu/_1463_ ( .A1(\mylsu/_0536_ ), .A2(\mylsu/_0584_ ), .A3(\mylsu/_0919_ ), .A4(\mylsu/_0535_ ), .ZN(\mylsu/_0299_ ) );
NAND3_X1 \mylsu/_1464_ ( .A1(\mylsu/_0584_ ), .A2(\mylsu/_0536_ ), .A3(\mylsu/_0535_ ), .ZN(\mylsu/_0300_ ) );
MUX2_X1 \mylsu/_1465_ ( .A(fanout_net_25 ), .B(\mylsu/_0266_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0234_ ) );
MUX2_X1 \mylsu/_1466_ ( .A(\mylsu/_0321_ ), .B(\mylsu/_0277_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0245_ ) );
MUX2_X1 \mylsu/_1467_ ( .A(\mylsu/_0332_ ), .B(\mylsu/_0288_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0256_ ) );
MUX2_X1 \mylsu/_1468_ ( .A(\mylsu/_0335_ ), .B(\mylsu/_0291_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0259_ ) );
MUX2_X1 \mylsu/_1469_ ( .A(\mylsu/_0336_ ), .B(\mylsu/_0292_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0260_ ) );
MUX2_X1 \mylsu/_1470_ ( .A(\mylsu/_0337_ ), .B(\mylsu/_0293_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0261_ ) );
MUX2_X1 \mylsu/_1471_ ( .A(\mylsu/_0338_ ), .B(\mylsu/_0294_ ), .S(\mylsu/_0578_ ), .Z(\mylsu/_0262_ ) );
BUF_X4 \mylsu/_1472_ ( .A(\mylsu/_0577_ ), .Z(\mylsu/_0585_ ) );
MUX2_X1 \mylsu/_1473_ ( .A(\mylsu/_0339_ ), .B(\mylsu/_0295_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0263_ ) );
MUX2_X1 \mylsu/_1474_ ( .A(\mylsu/_0340_ ), .B(\mylsu/_0296_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0264_ ) );
MUX2_X1 \mylsu/_1475_ ( .A(\mylsu/_0341_ ), .B(\mylsu/_0297_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0265_ ) );
MUX2_X1 \mylsu/_1476_ ( .A(\mylsu/_0311_ ), .B(\mylsu/_0267_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0235_ ) );
MUX2_X1 \mylsu/_1477_ ( .A(\mylsu/_0312_ ), .B(\mylsu/_0268_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0236_ ) );
MUX2_X1 \mylsu/_1478_ ( .A(\mylsu/_0313_ ), .B(\mylsu/_0269_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0237_ ) );
MUX2_X1 \mylsu/_1479_ ( .A(\mylsu/_0314_ ), .B(\mylsu/_0270_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0238_ ) );
MUX2_X1 \mylsu/_1480_ ( .A(\mylsu/_0315_ ), .B(\mylsu/_0271_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0239_ ) );
MUX2_X1 \mylsu/_1481_ ( .A(\mylsu/_0316_ ), .B(\mylsu/_0272_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0240_ ) );
MUX2_X1 \mylsu/_1482_ ( .A(\mylsu/_0317_ ), .B(\mylsu/_0273_ ), .S(\mylsu/_0585_ ), .Z(\mylsu/_0241_ ) );
BUF_X4 \mylsu/_1483_ ( .A(\mylsu/_0577_ ), .Z(\mylsu/_0586_ ) );
MUX2_X1 \mylsu/_1484_ ( .A(\mylsu/_0318_ ), .B(\mylsu/_0274_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0242_ ) );
MUX2_X1 \mylsu/_1485_ ( .A(\mylsu/_0319_ ), .B(\mylsu/_0275_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0243_ ) );
MUX2_X1 \mylsu/_1486_ ( .A(\mylsu/_0320_ ), .B(\mylsu/_0276_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0244_ ) );
MUX2_X1 \mylsu/_1487_ ( .A(\mylsu/_0322_ ), .B(\mylsu/_0278_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0246_ ) );
MUX2_X1 \mylsu/_1488_ ( .A(\mylsu/_0323_ ), .B(\mylsu/_0279_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0247_ ) );
MUX2_X1 \mylsu/_1489_ ( .A(\mylsu/_0324_ ), .B(\mylsu/_0280_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0248_ ) );
MUX2_X1 \mylsu/_1490_ ( .A(\mylsu/_0325_ ), .B(\mylsu/_0281_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0249_ ) );
MUX2_X1 \mylsu/_1491_ ( .A(\mylsu/_0326_ ), .B(\mylsu/_0282_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0250_ ) );
MUX2_X1 \mylsu/_1492_ ( .A(\mylsu/_0327_ ), .B(\mylsu/_0283_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0251_ ) );
MUX2_X1 \mylsu/_1493_ ( .A(\mylsu/_0328_ ), .B(\mylsu/_0284_ ), .S(\mylsu/_0586_ ), .Z(\mylsu/_0252_ ) );
MUX2_X1 \mylsu/_1494_ ( .A(\mylsu/_0329_ ), .B(\mylsu/_0285_ ), .S(\mylsu/_0577_ ), .Z(\mylsu/_0253_ ) );
MUX2_X1 \mylsu/_1495_ ( .A(\mylsu/_0330_ ), .B(\mylsu/_0286_ ), .S(\mylsu/_0577_ ), .Z(\mylsu/_0254_ ) );
MUX2_X1 \mylsu/_1496_ ( .A(\mylsu/_0331_ ), .B(\mylsu/_0287_ ), .S(\mylsu/_0577_ ), .Z(\mylsu/_0255_ ) );
MUX2_X1 \mylsu/_1497_ ( .A(\mylsu/_0333_ ), .B(\mylsu/_0289_ ), .S(\mylsu/_0577_ ), .Z(\mylsu/_0257_ ) );
MUX2_X1 \mylsu/_1498_ ( .A(\mylsu/_0334_ ), .B(\mylsu/_0290_ ), .S(\mylsu/_0577_ ), .Z(\mylsu/_0258_ ) );
INV_X1 \mylsu/_1499_ ( .A(\mylsu/_0839_ ), .ZN(\mylsu/_0587_ ) );
NOR3_X1 \mylsu/_1500_ ( .A1(\mylsu/_0587_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0947_ ) );
INV_X1 \mylsu/_1501_ ( .A(\mylsu/_0850_ ), .ZN(\mylsu/_0588_ ) );
NOR3_X1 \mylsu/_1502_ ( .A1(\mylsu/_0588_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0958_ ) );
INV_X1 \mylsu/_1503_ ( .A(\mylsu/_0861_ ), .ZN(\mylsu/_0589_ ) );
NOR3_X1 \mylsu/_1504_ ( .A1(\mylsu/_0589_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0969_ ) );
INV_X1 \mylsu/_1505_ ( .A(\mylsu/_0864_ ), .ZN(\mylsu/_0590_ ) );
NOR3_X1 \mylsu/_1506_ ( .A1(\mylsu/_0590_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0972_ ) );
INV_X1 \mylsu/_1507_ ( .A(\mylsu/_0865_ ), .ZN(\mylsu/_0591_ ) );
NOR3_X1 \mylsu/_1508_ ( .A1(\mylsu/_0591_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0973_ ) );
INV_X1 \mylsu/_1509_ ( .A(\mylsu/_0866_ ), .ZN(\mylsu/_0592_ ) );
NOR3_X1 \mylsu/_1510_ ( .A1(\mylsu/_0592_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0974_ ) );
INV_X1 \mylsu/_1511_ ( .A(\mylsu/_0867_ ), .ZN(\mylsu/_0593_ ) );
NOR3_X1 \mylsu/_1512_ ( .A1(\mylsu/_0593_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0975_ ) );
INV_X1 \mylsu/_1513_ ( .A(\mylsu/_0868_ ), .ZN(\mylsu/_0594_ ) );
NOR3_X1 \mylsu/_1514_ ( .A1(\mylsu/_0594_ ), .A2(fanout_net_25 ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_0976_ ) );
MUX2_X1 \mylsu/_1515_ ( .A(\mylsu/_0869_ ), .B(\mylsu/_0839_ ), .S(fanout_net_25 ), .Z(\mylsu/_0595_ ) );
INV_X2 \mylsu/_1516_ ( .A(\mylsu/_0321_ ), .ZN(\mylsu/_0596_ ) );
CLKBUF_X2 \mylsu/_1517_ ( .A(\mylsu/_0596_ ), .Z(\mylsu/_0597_ ) );
AND2_X1 \mylsu/_1518_ ( .A1(\mylsu/_0595_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0977_ ) );
MUX2_X1 \mylsu/_1519_ ( .A(\mylsu/_0870_ ), .B(\mylsu/_0850_ ), .S(fanout_net_25 ), .Z(\mylsu/_0598_ ) );
AND2_X1 \mylsu/_1520_ ( .A1(\mylsu/_0598_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0978_ ) );
MUX2_X1 \mylsu/_1521_ ( .A(\mylsu/_0840_ ), .B(\mylsu/_0861_ ), .S(fanout_net_25 ), .Z(\mylsu/_0599_ ) );
AND2_X1 \mylsu/_1522_ ( .A1(\mylsu/_0599_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0948_ ) );
MUX2_X1 \mylsu/_1523_ ( .A(\mylsu/_0841_ ), .B(\mylsu/_0864_ ), .S(fanout_net_25 ), .Z(\mylsu/_0600_ ) );
AND2_X1 \mylsu/_1524_ ( .A1(\mylsu/_0600_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0949_ ) );
MUX2_X1 \mylsu/_1525_ ( .A(\mylsu/_0842_ ), .B(\mylsu/_0865_ ), .S(fanout_net_25 ), .Z(\mylsu/_0601_ ) );
AND2_X1 \mylsu/_1526_ ( .A1(\mylsu/_0601_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0950_ ) );
MUX2_X1 \mylsu/_1527_ ( .A(\mylsu/_0843_ ), .B(\mylsu/_0866_ ), .S(fanout_net_25 ), .Z(\mylsu/_0602_ ) );
AND2_X1 \mylsu/_1528_ ( .A1(\mylsu/_0602_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0951_ ) );
MUX2_X1 \mylsu/_1529_ ( .A(\mylsu/_0844_ ), .B(\mylsu/_0867_ ), .S(fanout_net_25 ), .Z(\mylsu/_0603_ ) );
AND2_X1 \mylsu/_1530_ ( .A1(\mylsu/_0603_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0952_ ) );
MUX2_X1 \mylsu/_1531_ ( .A(\mylsu/_0845_ ), .B(\mylsu/_0868_ ), .S(fanout_net_25 ), .Z(\mylsu/_0604_ ) );
AND2_X1 \mylsu/_1532_ ( .A1(\mylsu/_0604_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_0953_ ) );
NOR2_X1 \mylsu/_1533_ ( .A1(\mylsu/_0587_ ), .A2(fanout_net_25 ), .ZN(\mylsu/_0605_ ) );
MUX2_X1 \mylsu/_1534_ ( .A(\mylsu/_0846_ ), .B(\mylsu/_0869_ ), .S(fanout_net_25 ), .Z(\mylsu/_0606_ ) );
MUX2_X1 \mylsu/_1535_ ( .A(\mylsu/_0605_ ), .B(\mylsu/_0606_ ), .S(\mylsu/_0597_ ), .Z(\mylsu/_0954_ ) );
NOR2_X1 \mylsu/_1536_ ( .A1(\mylsu/_0588_ ), .A2(fanout_net_25 ), .ZN(\mylsu/_0607_ ) );
MUX2_X1 \mylsu/_1537_ ( .A(\mylsu/_0847_ ), .B(\mylsu/_0870_ ), .S(fanout_net_25 ), .Z(\mylsu/_0608_ ) );
MUX2_X1 \mylsu/_1538_ ( .A(\mylsu/_0607_ ), .B(\mylsu/_0608_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0955_ ) );
NOR2_X1 \mylsu/_1539_ ( .A1(\mylsu/_0589_ ), .A2(fanout_net_25 ), .ZN(\mylsu/_0609_ ) );
MUX2_X1 \mylsu/_1540_ ( .A(\mylsu/_0848_ ), .B(\mylsu/_0840_ ), .S(fanout_net_25 ), .Z(\mylsu/_0610_ ) );
MUX2_X1 \mylsu/_1541_ ( .A(\mylsu/_0609_ ), .B(\mylsu/_0610_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0956_ ) );
NOR2_X1 \mylsu/_1542_ ( .A1(\mylsu/_0590_ ), .A2(fanout_net_25 ), .ZN(\mylsu/_0611_ ) );
MUX2_X1 \mylsu/_1543_ ( .A(\mylsu/_0849_ ), .B(\mylsu/_0841_ ), .S(fanout_net_25 ), .Z(\mylsu/_0612_ ) );
MUX2_X1 \mylsu/_1544_ ( .A(\mylsu/_0611_ ), .B(\mylsu/_0612_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0957_ ) );
NOR2_X1 \mylsu/_1545_ ( .A1(\mylsu/_0591_ ), .A2(fanout_net_25 ), .ZN(\mylsu/_0613_ ) );
MUX2_X1 \mylsu/_1546_ ( .A(\mylsu/_0851_ ), .B(\mylsu/_0842_ ), .S(fanout_net_25 ), .Z(\mylsu/_0614_ ) );
MUX2_X1 \mylsu/_1547_ ( .A(\mylsu/_0613_ ), .B(\mylsu/_0614_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0959_ ) );
NOR2_X1 \mylsu/_1548_ ( .A1(\mylsu/_0592_ ), .A2(fanout_net_25 ), .ZN(\mylsu/_0615_ ) );
MUX2_X1 \mylsu/_1549_ ( .A(\mylsu/_0852_ ), .B(\mylsu/_0843_ ), .S(fanout_net_25 ), .Z(\mylsu/_0616_ ) );
MUX2_X1 \mylsu/_1550_ ( .A(\mylsu/_0615_ ), .B(\mylsu/_0616_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0960_ ) );
NOR2_X1 \mylsu/_1551_ ( .A1(\mylsu/_0593_ ), .A2(\mylsu/_0310_ ), .ZN(\mylsu/_0617_ ) );
MUX2_X1 \mylsu/_1552_ ( .A(\mylsu/_0853_ ), .B(\mylsu/_0844_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0618_ ) );
MUX2_X1 \mylsu/_1553_ ( .A(\mylsu/_0617_ ), .B(\mylsu/_0618_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0961_ ) );
NOR2_X1 \mylsu/_1554_ ( .A1(\mylsu/_0594_ ), .A2(\mylsu/_0310_ ), .ZN(\mylsu/_0619_ ) );
MUX2_X1 \mylsu/_1555_ ( .A(\mylsu/_0854_ ), .B(\mylsu/_0845_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0620_ ) );
MUX2_X1 \mylsu/_1556_ ( .A(\mylsu/_0619_ ), .B(\mylsu/_0620_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_0962_ ) );
MUX2_X1 \mylsu/_1557_ ( .A(\mylsu/_0855_ ), .B(\mylsu/_0846_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0621_ ) );
MUX2_X1 \mylsu/_1558_ ( .A(\mylsu/_0621_ ), .B(\mylsu/_0595_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0963_ ) );
MUX2_X1 \mylsu/_1559_ ( .A(\mylsu/_0856_ ), .B(\mylsu/_0847_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0622_ ) );
MUX2_X1 \mylsu/_1560_ ( .A(\mylsu/_0622_ ), .B(\mylsu/_0598_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0964_ ) );
MUX2_X1 \mylsu/_1561_ ( .A(\mylsu/_0857_ ), .B(\mylsu/_0848_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0623_ ) );
MUX2_X1 \mylsu/_1562_ ( .A(\mylsu/_0623_ ), .B(\mylsu/_0599_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0965_ ) );
MUX2_X1 \mylsu/_1563_ ( .A(\mylsu/_0858_ ), .B(\mylsu/_0849_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0624_ ) );
MUX2_X1 \mylsu/_1564_ ( .A(\mylsu/_0624_ ), .B(\mylsu/_0600_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0966_ ) );
MUX2_X1 \mylsu/_1565_ ( .A(\mylsu/_0859_ ), .B(\mylsu/_0851_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0625_ ) );
MUX2_X1 \mylsu/_1566_ ( .A(\mylsu/_0625_ ), .B(\mylsu/_0601_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0967_ ) );
MUX2_X1 \mylsu/_1567_ ( .A(\mylsu/_0860_ ), .B(\mylsu/_0852_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0626_ ) );
MUX2_X1 \mylsu/_1568_ ( .A(\mylsu/_0626_ ), .B(\mylsu/_0602_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0968_ ) );
MUX2_X1 \mylsu/_1569_ ( .A(\mylsu/_0862_ ), .B(\mylsu/_0853_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0627_ ) );
MUX2_X1 \mylsu/_1570_ ( .A(\mylsu/_0627_ ), .B(\mylsu/_0603_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0970_ ) );
MUX2_X1 \mylsu/_1571_ ( .A(\mylsu/_0863_ ), .B(\mylsu/_0854_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0628_ ) );
MUX2_X1 \mylsu/_1572_ ( .A(\mylsu/_0628_ ), .B(\mylsu/_0604_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_0971_ ) );
NOR3_X1 \mylsu/_1573_ ( .A1(\mylsu/_0583_ ), .A2(\mylsu/_0310_ ), .A3(\mylsu/_0321_ ), .ZN(\mylsu/_1048_ ) );
MUX2_X1 \mylsu/_1574_ ( .A(\mylsu/_0919_ ), .B(\mylsu/_0918_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0629_ ) );
AND2_X1 \mylsu/_1575_ ( .A1(\mylsu/_0629_ ), .A2(\mylsu/_0597_ ), .ZN(\mylsu/_1049_ ) );
NOR2_X1 \mylsu/_1576_ ( .A1(\mylsu/_0583_ ), .A2(\mylsu/_0310_ ), .ZN(\mylsu/_0630_ ) );
MUX2_X1 \mylsu/_1577_ ( .A(\mylsu/_0920_ ), .B(\mylsu/_0919_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0631_ ) );
MUX2_X1 \mylsu/_1578_ ( .A(\mylsu/_0630_ ), .B(\mylsu/_0631_ ), .S(\mylsu/_0596_ ), .Z(\mylsu/_1050_ ) );
MUX2_X1 \mylsu/_1579_ ( .A(\mylsu/_0921_ ), .B(\mylsu/_0920_ ), .S(\mylsu/_0310_ ), .Z(\mylsu/_0632_ ) );
MUX2_X1 \mylsu/_1580_ ( .A(\mylsu/_0632_ ), .B(\mylsu/_0629_ ), .S(\mylsu/_0321_ ), .Z(\mylsu/_1051_ ) );
BUF_X4 \mylsu/_1581_ ( .A(\mylsu/_0567_ ), .Z(\mylsu/_0633_ ) );
MUX2_X1 \mylsu/_1582_ ( .A(\mylsu/_0942_ ), .B(\mylsu/_0342_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0081_ ) );
MUX2_X1 \mylsu/_1583_ ( .A(\mylsu/_0943_ ), .B(\mylsu/_0343_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0082_ ) );
MUX2_X1 \mylsu/_1584_ ( .A(\mylsu/_0944_ ), .B(\mylsu/_0344_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0083_ ) );
MUX2_X1 \mylsu/_1585_ ( .A(\mylsu/_0945_ ), .B(\mylsu/_0345_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0084_ ) );
MUX2_X1 \mylsu/_1586_ ( .A(\mylsu/_0946_ ), .B(\mylsu/_0346_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0085_ ) );
NOR2_X1 \mylsu/_1587_ ( .A1(\mylsu/_0923_ ), .A2(\mylsu/_0924_ ), .ZN(\mylsu/_0634_ ) );
NOR2_X4 \mylsu/_1588_ ( .A1(\mylsu/_0550_ ), .A2(\mylsu/_0634_ ), .ZN(\mylsu/_0635_ ) );
AND2_X1 \mylsu/_1589_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0551_ ), .ZN(\mylsu/_0636_ ) );
INV_X1 \mylsu/_1590_ ( .A(\mylsu/_0636_ ), .ZN(\mylsu/_0637_ ) );
AOI21_X1 \mylsu/_1591_ ( .A(\mylsu/_0930_ ), .B1(\mylsu/_0637_ ), .B2(\mylsu/_0633_ ), .ZN(\mylsu/_0638_ ) );
NAND2_X1 \mylsu/_1592_ ( .A1(\mylsu/_0534_ ), .A2(\mylsu/_0925_ ), .ZN(\mylsu/_0639_ ) );
AND2_X1 \mylsu/_1593_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0639_ ), .ZN(\mylsu/_0640_ ) );
BUF_X4 \mylsu/_1594_ ( .A(\mylsu/_0640_ ), .Z(\mylsu/_0641_ ) );
BUF_X8 \mylsu/_1595_ ( .A(\mylsu/_0641_ ), .Z(\mylsu/_0642_ ) );
AND2_X1 \mylsu/_1596_ ( .A1(\mylsu/_0637_ ), .A2(\mylsu/_0642_ ), .ZN(\mylsu/_0643_ ) );
INV_X1 \mylsu/_1597_ ( .A(\mylsu/_0549_ ), .ZN(\mylsu/_0644_ ) );
NOR3_X1 \mylsu/_1598_ ( .A1(\mylsu/_0644_ ), .A2(fanout_net_26 ), .A3(\mylsu/_0310_ ), .ZN(\mylsu/_0645_ ) );
AOI21_X1 \mylsu/_1599_ ( .A(\mylsu/_0638_ ), .B1(\mylsu/_0643_ ), .B2(\mylsu/_0645_ ), .ZN(\mylsu/_0086_ ) );
BUF_X2 \mylsu/_1600_ ( .A(\mylsu/_0635_ ), .Z(\mylsu/_0646_ ) );
CLKBUF_X2 \mylsu/_1601_ ( .A(\mylsu/_0639_ ), .Z(\mylsu/_0647_ ) );
AND3_X1 \mylsu/_1602_ ( .A1(\mylsu/_0646_ ), .A2(\mylsu/_0321_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0648_ ) );
INV_X1 \mylsu/_1603_ ( .A(\mylsu/_0567_ ), .ZN(\mylsu/_0649_ ) );
NOR2_X2 \mylsu/_1604_ ( .A1(\mylsu/_0636_ ), .A2(\mylsu/_0649_ ), .ZN(\mylsu/_0650_ ) );
BUF_X4 \mylsu/_1605_ ( .A(\mylsu/_0650_ ), .Z(\mylsu/_0651_ ) );
MUX2_X1 \mylsu/_1606_ ( .A(\mylsu/_0933_ ), .B(\mylsu/_0648_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0087_ ) );
AND3_X1 \mylsu/_1607_ ( .A1(\mylsu/_0646_ ), .A2(\mylsu/_0332_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0652_ ) );
MUX2_X1 \mylsu/_1608_ ( .A(\mylsu/_0934_ ), .B(\mylsu/_0652_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0088_ ) );
AND3_X1 \mylsu/_1609_ ( .A1(\mylsu/_0646_ ), .A2(\mylsu/_0335_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0653_ ) );
MUX2_X1 \mylsu/_1610_ ( .A(\mylsu/_0935_ ), .B(\mylsu/_0653_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0089_ ) );
AND3_X1 \mylsu/_1611_ ( .A1(\mylsu/_0646_ ), .A2(\mylsu/_0336_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0654_ ) );
MUX2_X1 \mylsu/_1612_ ( .A(\mylsu/_0936_ ), .B(\mylsu/_0654_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0090_ ) );
AND3_X1 \mylsu/_1613_ ( .A1(\mylsu/_0646_ ), .A2(\mylsu/_0337_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0655_ ) );
MUX2_X1 \mylsu/_1614_ ( .A(\mylsu/_0937_ ), .B(\mylsu/_0655_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0091_ ) );
NAND3_X1 \mylsu/_1615_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0338_ ), .A3(\mylsu/_0639_ ), .ZN(\mylsu/_0656_ ) );
NAND3_X1 \mylsu/_1616_ ( .A1(\mylsu/_0656_ ), .A2(\mylsu/_0646_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0657_ ) );
MUX2_X1 \mylsu/_1617_ ( .A(\mylsu/_0938_ ), .B(\mylsu/_0657_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0092_ ) );
AND3_X1 \mylsu/_1618_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0339_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0658_ ) );
MUX2_X1 \mylsu/_1619_ ( .A(\mylsu/_0939_ ), .B(\mylsu/_0658_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0093_ ) );
NAND3_X1 \mylsu/_1620_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0340_ ), .A3(\mylsu/_0639_ ), .ZN(\mylsu/_0659_ ) );
NAND3_X1 \mylsu/_1621_ ( .A1(\mylsu/_0659_ ), .A2(\mylsu/_0646_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0660_ ) );
MUX2_X1 \mylsu/_1622_ ( .A(\mylsu/_0940_ ), .B(\mylsu/_0660_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0094_ ) );
NAND3_X1 \mylsu/_1623_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0341_ ), .A3(\mylsu/_0639_ ), .ZN(\mylsu/_0661_ ) );
NAND3_X1 \mylsu/_1624_ ( .A1(\mylsu/_0661_ ), .A2(\mylsu/_0646_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0662_ ) );
MUX2_X1 \mylsu/_1625_ ( .A(\mylsu/_0941_ ), .B(\mylsu/_0662_ ), .S(\mylsu/_0651_ ), .Z(\mylsu/_0095_ ) );
AND3_X1 \mylsu/_1626_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0311_ ), .A3(\mylsu/_0639_ ), .ZN(\mylsu/_0663_ ) );
BUF_X4 \mylsu/_1627_ ( .A(\mylsu/_0650_ ), .Z(\mylsu/_0664_ ) );
MUX2_X1 \mylsu/_1628_ ( .A(\mylsu/_0931_ ), .B(\mylsu/_0663_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0096_ ) );
AND3_X1 \mylsu/_1629_ ( .A1(\mylsu/_0635_ ), .A2(\mylsu/_0312_ ), .A3(\mylsu/_0639_ ), .ZN(\mylsu/_0665_ ) );
MUX2_X1 \mylsu/_1630_ ( .A(\mylsu/_0932_ ), .B(\mylsu/_0665_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0097_ ) );
NOR2_X1 \mylsu/_1631_ ( .A1(\mylsu/_0547_ ), .A2(\mylsu/_0913_ ), .ZN(\mylsu/_0666_ ) );
OAI21_X4 \mylsu/_1632_ ( .A(\mylsu/_0548_ ), .B1(\mylsu/_0549_ ), .B2(\mylsu/_0666_ ), .ZN(\mylsu/_0667_ ) );
BUF_X4 \mylsu/_1633_ ( .A(\mylsu/_0667_ ), .Z(\mylsu/_0668_ ) );
OAI21_X1 \mylsu/_1634_ ( .A(\mylsu/_1011_ ), .B1(\mylsu/_0668_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0669_ ) );
INV_X32 \mylsu/_1635_ ( .A(\mylsu/_0046_ ), .ZN(\mylsu/_0670_ ) );
NOR2_X1 \mylsu/_1636_ ( .A1(\mylsu/_0670_ ), .A2(\mylsu/_0057_ ), .ZN(\mylsu/_0671_ ) );
INV_X2 \mylsu/_1637_ ( .A(\mylsu/_0671_ ), .ZN(\mylsu/_0672_ ) );
INV_X8 \mylsu/_1638_ ( .A(\mylsu/_0057_ ), .ZN(\mylsu/_0673_ ) );
NOR2_X4 \mylsu/_1639_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .ZN(\mylsu/_0674_ ) );
INV_X1 \mylsu/_1640_ ( .A(\mylsu/_0822_ ), .ZN(\mylsu/_0675_ ) );
OAI21_X1 \mylsu/_1641_ ( .A(\mylsu/_0672_ ), .B1(\mylsu/_0674_ ), .B2(\mylsu/_0675_ ), .ZN(\mylsu/_0676_ ) );
NOR2_X4 \mylsu/_1642_ ( .A1(\mylsu/_0927_ ), .A2(\mylsu/_0926_ ), .ZN(\mylsu/_0677_ ) );
AND2_X1 \mylsu/_1643_ ( .A1(\mylsu/_0677_ ), .A2(\mylsu/_0013_ ), .ZN(\mylsu/_0678_ ) );
BUF_X2 \mylsu/_1644_ ( .A(\mylsu/_0678_ ), .Z(\mylsu/_0679_ ) );
NAND2_X1 \mylsu/_1645_ ( .A1(\mylsu/_0926_ ), .A2(\mylsu/_0013_ ), .ZN(\mylsu/_0680_ ) );
NOR2_X2 \mylsu/_1646_ ( .A1(\mylsu/_0680_ ), .A2(\mylsu/_0927_ ), .ZN(\mylsu/_0681_ ) );
OAI221_X1 \mylsu/_1647_ ( .A(\mylsu/_0676_ ), .B1(\mylsu/_0836_ ), .B2(\mylsu/_0672_ ), .C1(\mylsu/_0679_ ), .C2(\mylsu/_0681_ ), .ZN(\mylsu/_0682_ ) );
NOR2_X4 \mylsu/_1648_ ( .A1(\mylsu/_0679_ ), .A2(\mylsu/_0681_ ), .ZN(\mylsu/_0683_ ) );
BUF_X4 \mylsu/_1649_ ( .A(\mylsu/_0683_ ), .Z(\mylsu/_0684_ ) );
OAI21_X1 \mylsu/_1650_ ( .A(\mylsu/_0813_ ), .B1(\mylsu/_0684_ ), .B2(\mylsu/_0674_ ), .ZN(\mylsu/_0685_ ) );
NAND2_X4 \mylsu/_1651_ ( .A1(\mylsu/_0927_ ), .A2(\mylsu/_0013_ ), .ZN(\mylsu/_0686_ ) );
NOR2_X1 \mylsu/_1652_ ( .A1(\mylsu/_0686_ ), .A2(\mylsu/_0926_ ), .ZN(\mylsu/_0687_ ) );
NAND2_X1 \mylsu/_1653_ ( .A1(\mylsu/_0927_ ), .A2(\mylsu/_0926_ ), .ZN(\mylsu/_0688_ ) );
NOR2_X2 \mylsu/_1654_ ( .A1(\mylsu/_0688_ ), .A2(\mylsu/_0928_ ), .ZN(\mylsu/_0689_ ) );
NOR2_X2 \mylsu/_1655_ ( .A1(\mylsu/_0687_ ), .A2(\mylsu/_0689_ ), .ZN(\mylsu/_0690_ ) );
AND2_X1 \mylsu/_1656_ ( .A1(\mylsu/_0683_ ), .A2(\mylsu/_0690_ ), .ZN(\mylsu/_0691_ ) );
OAI21_X1 \mylsu/_1657_ ( .A(\mylsu/_0682_ ), .B1(\mylsu/_0685_ ), .B2(\mylsu/_0691_ ), .ZN(\mylsu/_0692_ ) );
NOR2_X4 \mylsu/_1658_ ( .A1(\mylsu/_0046_ ), .A2(\mylsu/_0057_ ), .ZN(\mylsu/_0693_ ) );
INV_X4 \mylsu/_1659_ ( .A(\mylsu/_0693_ ), .ZN(\mylsu/_0694_ ) );
NAND2_X1 \mylsu/_1660_ ( .A1(\mylsu/_0692_ ), .A2(\mylsu/_0694_ ), .ZN(\mylsu/_0695_ ) );
BUF_X4 \mylsu/_1661_ ( .A(\mylsu/_0693_ ), .Z(\mylsu/_0696_ ) );
OAI21_X1 \mylsu/_1662_ ( .A(\mylsu/_0806_ ), .B1(\mylsu/_0691_ ), .B2(\mylsu/_0696_ ), .ZN(\mylsu/_0697_ ) );
AND3_X1 \mylsu/_1663_ ( .A1(\mylsu/_0695_ ), .A2(fanout_net_27 ), .A3(\mylsu/_0697_ ), .ZN(\mylsu/_0698_ ) );
NOR2_X4 \mylsu/_1664_ ( .A1(\mylsu/_0667_ ), .A2(fanout_net_26 ), .ZN(\mylsu/_0699_ ) );
BUF_X4 \mylsu/_1665_ ( .A(\mylsu/_0699_ ), .Z(\mylsu/_0700_ ) );
OAI21_X1 \mylsu/_1666_ ( .A(\mylsu/_0700_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0871_ ), .ZN(\mylsu/_0701_ ) );
OAI21_X1 \mylsu/_1667_ ( .A(\mylsu/_0669_ ), .B1(\mylsu/_0698_ ), .B2(\mylsu/_0701_ ), .ZN(\mylsu/_0098_ ) );
OAI21_X1 \mylsu/_1668_ ( .A(\mylsu/_1022_ ), .B1(\mylsu/_0668_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0702_ ) );
AND3_X1 \mylsu/_1669_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .A3(\mylsu/_0837_ ), .ZN(\mylsu/_0703_ ) );
MUX2_X1 \mylsu/_1670_ ( .A(\mylsu/_0823_ ), .B(\mylsu/_0814_ ), .S(\mylsu/_0674_ ), .Z(\mylsu/_0704_ ) );
AOI211_X4 \mylsu/_1671_ ( .A(\mylsu/_0683_ ), .B(\mylsu/_0703_ ), .C1(\mylsu/_0704_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0705_ ) );
BUF_X4 \mylsu/_1672_ ( .A(\mylsu/_0690_ ), .Z(\mylsu/_0706_ ) );
NOR4_X1 \mylsu/_1673_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0679_ ), .A3(\mylsu/_0814_ ), .A4(\mylsu/_0681_ ), .ZN(\mylsu/_0707_ ) );
OAI21_X1 \mylsu/_1674_ ( .A(\mylsu/_0694_ ), .B1(\mylsu/_0705_ ), .B2(\mylsu/_0707_ ), .ZN(\mylsu/_0708_ ) );
NOR2_X1 \mylsu/_1675_ ( .A1(\mylsu/_0691_ ), .A2(\mylsu/_0696_ ), .ZN(\mylsu/_0709_ ) );
OR2_X1 \mylsu/_1676_ ( .A1(\mylsu/_0709_ ), .A2(\mylsu/_0817_ ), .ZN(\mylsu/_0710_ ) );
AOI21_X1 \mylsu/_1677_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0708_ ), .B2(\mylsu/_0710_ ), .ZN(\mylsu/_0711_ ) );
OAI21_X1 \mylsu/_1678_ ( .A(\mylsu/_0700_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0882_ ), .ZN(\mylsu/_0712_ ) );
OAI21_X1 \mylsu/_1679_ ( .A(\mylsu/_0702_ ), .B1(\mylsu/_0711_ ), .B2(\mylsu/_0712_ ), .ZN(\mylsu/_0099_ ) );
OAI21_X1 \mylsu/_1680_ ( .A(\mylsu/_1033_ ), .B1(\mylsu/_0668_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0713_ ) );
AND3_X1 \mylsu/_1681_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .A3(\mylsu/_0807_ ), .ZN(\mylsu/_0714_ ) );
MUX2_X1 \mylsu/_1682_ ( .A(\mylsu/_0824_ ), .B(\mylsu/_0815_ ), .S(\mylsu/_0674_ ), .Z(\mylsu/_0715_ ) );
AOI211_X4 \mylsu/_1683_ ( .A(\mylsu/_0683_ ), .B(\mylsu/_0714_ ), .C1(\mylsu/_0715_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0716_ ) );
NOR4_X1 \mylsu/_1684_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0679_ ), .A3(\mylsu/_0815_ ), .A4(\mylsu/_0681_ ), .ZN(\mylsu/_0717_ ) );
OAI21_X1 \mylsu/_1685_ ( .A(\mylsu/_0694_ ), .B1(\mylsu/_0716_ ), .B2(\mylsu/_0717_ ), .ZN(\mylsu/_0718_ ) );
OR2_X1 \mylsu/_1686_ ( .A1(\mylsu/_0709_ ), .A2(\mylsu/_0828_ ), .ZN(\mylsu/_0719_ ) );
AOI21_X1 \mylsu/_1687_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0718_ ), .B2(\mylsu/_0719_ ), .ZN(\mylsu/_0720_ ) );
OAI21_X1 \mylsu/_1688_ ( .A(\mylsu/_0700_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0893_ ), .ZN(\mylsu/_0721_ ) );
OAI21_X1 \mylsu/_1689_ ( .A(\mylsu/_0713_ ), .B1(\mylsu/_0720_ ), .B2(\mylsu/_0721_ ), .ZN(\mylsu/_0100_ ) );
OAI21_X1 \mylsu/_1690_ ( .A(\mylsu/_1036_ ), .B1(\mylsu/_0668_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0722_ ) );
AND3_X1 \mylsu/_1691_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .A3(\mylsu/_0808_ ), .ZN(\mylsu/_0723_ ) );
MUX2_X1 \mylsu/_1692_ ( .A(\mylsu/_0825_ ), .B(\mylsu/_0816_ ), .S(\mylsu/_0674_ ), .Z(\mylsu/_0724_ ) );
AOI211_X4 \mylsu/_1693_ ( .A(\mylsu/_0683_ ), .B(\mylsu/_0723_ ), .C1(\mylsu/_0724_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0725_ ) );
NOR4_X1 \mylsu/_1694_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0679_ ), .A3(\mylsu/_0816_ ), .A4(\mylsu/_0681_ ), .ZN(\mylsu/_0726_ ) );
OAI21_X1 \mylsu/_1695_ ( .A(\mylsu/_0694_ ), .B1(\mylsu/_0725_ ), .B2(\mylsu/_0726_ ), .ZN(\mylsu/_0727_ ) );
OR2_X1 \mylsu/_1696_ ( .A1(\mylsu/_0709_ ), .A2(\mylsu/_0831_ ), .ZN(\mylsu/_0728_ ) );
AOI21_X1 \mylsu/_1697_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0727_ ), .B2(\mylsu/_0728_ ), .ZN(\mylsu/_0729_ ) );
OAI21_X1 \mylsu/_1698_ ( .A(\mylsu/_0700_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0896_ ), .ZN(\mylsu/_0730_ ) );
OAI21_X1 \mylsu/_1699_ ( .A(\mylsu/_0722_ ), .B1(\mylsu/_0729_ ), .B2(\mylsu/_0730_ ), .ZN(\mylsu/_0101_ ) );
OAI21_X1 \mylsu/_1700_ ( .A(\mylsu/_1037_ ), .B1(\mylsu/_0668_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0731_ ) );
AND3_X1 \mylsu/_1701_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .A3(\mylsu/_0809_ ), .ZN(\mylsu/_0732_ ) );
MUX2_X1 \mylsu/_1702_ ( .A(\mylsu/_0826_ ), .B(\mylsu/_0818_ ), .S(\mylsu/_0674_ ), .Z(\mylsu/_0733_ ) );
AOI211_X4 \mylsu/_1703_ ( .A(\mylsu/_0683_ ), .B(\mylsu/_0732_ ), .C1(\mylsu/_0733_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0734_ ) );
NOR4_X1 \mylsu/_1704_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0679_ ), .A3(\mylsu/_0818_ ), .A4(\mylsu/_0681_ ), .ZN(\mylsu/_0735_ ) );
OAI21_X1 \mylsu/_1705_ ( .A(\mylsu/_0694_ ), .B1(\mylsu/_0734_ ), .B2(\mylsu/_0735_ ), .ZN(\mylsu/_0736_ ) );
OR2_X1 \mylsu/_1706_ ( .A1(\mylsu/_0709_ ), .A2(\mylsu/_0832_ ), .ZN(\mylsu/_0737_ ) );
AOI21_X1 \mylsu/_1707_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0736_ ), .B2(\mylsu/_0737_ ), .ZN(\mylsu/_0738_ ) );
OAI21_X1 \mylsu/_1708_ ( .A(\mylsu/_0700_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0897_ ), .ZN(\mylsu/_0739_ ) );
OAI21_X1 \mylsu/_1709_ ( .A(\mylsu/_0731_ ), .B1(\mylsu/_0738_ ), .B2(\mylsu/_0739_ ), .ZN(\mylsu/_0102_ ) );
OAI21_X1 \mylsu/_1710_ ( .A(\mylsu/_1038_ ), .B1(\mylsu/_0667_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0740_ ) );
AND3_X1 \mylsu/_1711_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .A3(\mylsu/_0810_ ), .ZN(\mylsu/_0741_ ) );
MUX2_X1 \mylsu/_1712_ ( .A(\mylsu/_0827_ ), .B(\mylsu/_0819_ ), .S(\mylsu/_0674_ ), .Z(\mylsu/_0742_ ) );
AOI211_X4 \mylsu/_1713_ ( .A(\mylsu/_0683_ ), .B(\mylsu/_0741_ ), .C1(\mylsu/_0742_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0743_ ) );
NOR4_X1 \mylsu/_1714_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0679_ ), .A3(\mylsu/_0819_ ), .A4(\mylsu/_0681_ ), .ZN(\mylsu/_0744_ ) );
OAI21_X1 \mylsu/_1715_ ( .A(\mylsu/_0694_ ), .B1(\mylsu/_0743_ ), .B2(\mylsu/_0744_ ), .ZN(\mylsu/_0745_ ) );
OR2_X1 \mylsu/_1716_ ( .A1(\mylsu/_0709_ ), .A2(\mylsu/_0833_ ), .ZN(\mylsu/_0746_ ) );
AOI21_X1 \mylsu/_1717_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0745_ ), .B2(\mylsu/_0746_ ), .ZN(\mylsu/_0747_ ) );
OAI21_X1 \mylsu/_1718_ ( .A(\mylsu/_0699_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0898_ ), .ZN(\mylsu/_0748_ ) );
OAI21_X1 \mylsu/_1719_ ( .A(\mylsu/_0740_ ), .B1(\mylsu/_0747_ ), .B2(\mylsu/_0748_ ), .ZN(\mylsu/_0103_ ) );
OAI21_X1 \mylsu/_1720_ ( .A(\mylsu/_1039_ ), .B1(\mylsu/_0667_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0749_ ) );
AND3_X1 \mylsu/_1721_ ( .A1(\mylsu/_0673_ ), .A2(\mylsu/_0046_ ), .A3(\mylsu/_0811_ ), .ZN(\mylsu/_0750_ ) );
MUX2_X1 \mylsu/_1722_ ( .A(\mylsu/_0829_ ), .B(\mylsu/_0820_ ), .S(\mylsu/_0674_ ), .Z(\mylsu/_0751_ ) );
AOI211_X4 \mylsu/_1723_ ( .A(\mylsu/_0683_ ), .B(\mylsu/_0750_ ), .C1(\mylsu/_0751_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0752_ ) );
NOR4_X1 \mylsu/_1724_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0679_ ), .A3(\mylsu/_0820_ ), .A4(\mylsu/_0681_ ), .ZN(\mylsu/_0753_ ) );
OAI21_X1 \mylsu/_1725_ ( .A(\mylsu/_0694_ ), .B1(\mylsu/_0752_ ), .B2(\mylsu/_0753_ ), .ZN(\mylsu/_0754_ ) );
OR2_X1 \mylsu/_1726_ ( .A1(\mylsu/_0709_ ), .A2(\mylsu/_0834_ ), .ZN(\mylsu/_0755_ ) );
AOI21_X1 \mylsu/_1727_ ( .A(\mylsu/_0575_ ), .B1(\mylsu/_0754_ ), .B2(\mylsu/_0755_ ), .ZN(\mylsu/_0756_ ) );
OAI21_X1 \mylsu/_1728_ ( .A(\mylsu/_0699_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0899_ ), .ZN(\mylsu/_0757_ ) );
OAI21_X1 \mylsu/_1729_ ( .A(\mylsu/_0749_ ), .B1(\mylsu/_0756_ ), .B2(\mylsu/_0757_ ), .ZN(\mylsu/_0104_ ) );
NOR2_X1 \mylsu/_1730_ ( .A1(\mylsu/_0700_ ), .A2(\mylsu/_1040_ ), .ZN(\mylsu/_0758_ ) );
AOI211_X2 \mylsu/_1731_ ( .A(fanout_net_26 ), .B(\mylsu/_0667_ ), .C1(\mylsu/_0575_ ), .C2(\mylsu/_0900_ ), .ZN(\mylsu/_0759_ ) );
NAND3_X1 \mylsu/_1732_ ( .A1(\mylsu/_0670_ ), .A2(\mylsu/_0057_ ), .A3(\mylsu/_0821_ ), .ZN(\mylsu/_0760_ ) );
INV_X1 \mylsu/_1733_ ( .A(\mylsu/_0830_ ), .ZN(\mylsu/_0761_ ) );
OAI211_X2 \mylsu/_1734_ ( .A(\mylsu/_0672_ ), .B(\mylsu/_0760_ ), .C1(\mylsu/_0761_ ), .C2(\mylsu/_0674_ ), .ZN(\mylsu/_0762_ ) );
OAI211_X2 \mylsu/_1735_ ( .A(\mylsu/_0762_ ), .B(\mylsu/_0694_ ), .C1(\mylsu/_0812_ ), .C2(\mylsu/_0672_ ), .ZN(\mylsu/_0763_ ) );
INV_X1 \mylsu/_1736_ ( .A(\mylsu/_0684_ ), .ZN(\mylsu/_0764_ ) );
NAND3_X1 \mylsu/_1737_ ( .A1(\mylsu/_0670_ ), .A2(\mylsu/_0673_ ), .A3(\mylsu/_0835_ ), .ZN(\mylsu/_0765_ ) );
NAND3_X1 \mylsu/_1738_ ( .A1(\mylsu/_0763_ ), .A2(\mylsu/_0764_ ), .A3(\mylsu/_0765_ ), .ZN(\mylsu/_0766_ ) );
INV_X1 \mylsu/_1739_ ( .A(\mylsu/_0821_ ), .ZN(\mylsu/_0767_ ) );
OR3_X1 \mylsu/_1740_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0767_ ), .A3(\mylsu/_0693_ ), .ZN(\mylsu/_0768_ ) );
OAI21_X1 \mylsu/_1741_ ( .A(\mylsu/_0835_ ), .B1(\mylsu/_0706_ ), .B2(\mylsu/_0696_ ), .ZN(\mylsu/_0769_ ) );
NAND3_X1 \mylsu/_1742_ ( .A1(\mylsu/_0768_ ), .A2(\mylsu/_0769_ ), .A3(\mylsu/_0684_ ), .ZN(\mylsu/_0770_ ) );
NAND3_X1 \mylsu/_1743_ ( .A1(\mylsu/_0766_ ), .A2(\mylsu/_0770_ ), .A3(fanout_net_27 ), .ZN(\mylsu/_0771_ ) );
AOI21_X1 \mylsu/_1744_ ( .A(\mylsu/_0758_ ), .B1(\mylsu/_0759_ ), .B2(\mylsu/_0771_ ), .ZN(\mylsu/_0105_ ) );
NAND2_X2 \mylsu/_1745_ ( .A1(\mylsu/_0763_ ), .A2(\mylsu/_0765_ ), .ZN(\mylsu/_0347_ ) );
AND2_X2 \mylsu/_1746_ ( .A1(\mylsu/_0347_ ), .A2(\mylsu/_0679_ ), .ZN(\mylsu/_0348_ ) );
NOR2_X4 \mylsu/_1747_ ( .A1(\mylsu/_0348_ ), .A2(\mylsu/_0547_ ), .ZN(\mylsu/_0349_ ) );
NOR3_X1 \mylsu/_1748_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0822_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0350_ ) );
NOR2_X4 \mylsu/_1749_ ( .A1(\mylsu/_0690_ ), .A2(\mylsu/_0693_ ), .ZN(\mylsu/_0351_ ) );
OAI21_X1 \mylsu/_1750_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0836_ ), .ZN(\mylsu/_0352_ ) );
OAI21_X1 \mylsu/_1751_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0350_ ), .B2(\mylsu/_0352_ ), .ZN(\mylsu/_0353_ ) );
BUF_X8 \mylsu/_1752_ ( .A(\mylsu/_0699_ ), .Z(\mylsu/_0354_ ) );
OAI211_X2 \mylsu/_1753_ ( .A(\mylsu/_0353_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0901_ ), .ZN(\mylsu/_0355_ ) );
BUF_X4 \mylsu/_1754_ ( .A(\mylsu/_0667_ ), .Z(\mylsu/_0356_ ) );
OAI21_X1 \mylsu/_1755_ ( .A(\mylsu/_1041_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0357_ ) );
NAND2_X1 \mylsu/_1756_ ( .A1(\mylsu/_0355_ ), .A2(\mylsu/_0357_ ), .ZN(\mylsu/_0106_ ) );
NOR3_X1 \mylsu/_1757_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0823_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0358_ ) );
OAI21_X1 \mylsu/_1758_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0837_ ), .ZN(\mylsu/_0359_ ) );
OAI21_X1 \mylsu/_1759_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0358_ ), .B2(\mylsu/_0359_ ), .ZN(\mylsu/_0360_ ) );
OAI211_X2 \mylsu/_1760_ ( .A(\mylsu/_0360_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0902_ ), .ZN(\mylsu/_0361_ ) );
OAI21_X1 \mylsu/_1761_ ( .A(\mylsu/_1042_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0362_ ) );
NAND2_X1 \mylsu/_1762_ ( .A1(\mylsu/_0361_ ), .A2(\mylsu/_0362_ ), .ZN(\mylsu/_0107_ ) );
NOR3_X1 \mylsu/_1763_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0824_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0363_ ) );
OAI21_X1 \mylsu/_1764_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0807_ ), .ZN(\mylsu/_0364_ ) );
OAI21_X1 \mylsu/_1765_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0363_ ), .B2(\mylsu/_0364_ ), .ZN(\mylsu/_0365_ ) );
OAI211_X2 \mylsu/_1766_ ( .A(\mylsu/_0365_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0872_ ), .ZN(\mylsu/_0366_ ) );
OAI21_X1 \mylsu/_1767_ ( .A(\mylsu/_1012_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0367_ ) );
NAND2_X1 \mylsu/_1768_ ( .A1(\mylsu/_0366_ ), .A2(\mylsu/_0367_ ), .ZN(\mylsu/_0108_ ) );
NOR3_X1 \mylsu/_1769_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0825_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0368_ ) );
OAI21_X1 \mylsu/_1770_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0808_ ), .ZN(\mylsu/_0369_ ) );
OAI21_X2 \mylsu/_1771_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0368_ ), .B2(\mylsu/_0369_ ), .ZN(\mylsu/_0370_ ) );
OAI211_X2 \mylsu/_1772_ ( .A(\mylsu/_0370_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0873_ ), .ZN(\mylsu/_0371_ ) );
OAI21_X1 \mylsu/_1773_ ( .A(\mylsu/_1013_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0372_ ) );
NAND2_X1 \mylsu/_1774_ ( .A1(\mylsu/_0371_ ), .A2(\mylsu/_0372_ ), .ZN(\mylsu/_0109_ ) );
NOR3_X1 \mylsu/_1775_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0826_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0373_ ) );
OAI21_X1 \mylsu/_1776_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0809_ ), .ZN(\mylsu/_0374_ ) );
OAI21_X1 \mylsu/_1777_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0373_ ), .B2(\mylsu/_0374_ ), .ZN(\mylsu/_0375_ ) );
OAI211_X2 \mylsu/_1778_ ( .A(\mylsu/_0375_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0874_ ), .ZN(\mylsu/_0376_ ) );
OAI21_X1 \mylsu/_1779_ ( .A(\mylsu/_1014_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0377_ ) );
NAND2_X1 \mylsu/_1780_ ( .A1(\mylsu/_0376_ ), .A2(\mylsu/_0377_ ), .ZN(\mylsu/_0110_ ) );
NOR3_X1 \mylsu/_1781_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0827_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0378_ ) );
OAI21_X1 \mylsu/_1782_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0810_ ), .ZN(\mylsu/_0379_ ) );
OAI21_X1 \mylsu/_1783_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0378_ ), .B2(\mylsu/_0379_ ), .ZN(\mylsu/_0380_ ) );
OAI211_X2 \mylsu/_1784_ ( .A(\mylsu/_0380_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0875_ ), .ZN(\mylsu/_0381_ ) );
OAI21_X1 \mylsu/_1785_ ( .A(\mylsu/_1015_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0382_ ) );
NAND2_X1 \mylsu/_1786_ ( .A1(\mylsu/_0381_ ), .A2(\mylsu/_0382_ ), .ZN(\mylsu/_0111_ ) );
NOR3_X1 \mylsu/_1787_ ( .A1(\mylsu/_0706_ ), .A2(\mylsu/_0829_ ), .A3(\mylsu/_0696_ ), .ZN(\mylsu/_0383_ ) );
OAI21_X1 \mylsu/_1788_ ( .A(\mylsu/_0684_ ), .B1(\mylsu/_0351_ ), .B2(\mylsu/_0811_ ), .ZN(\mylsu/_0384_ ) );
OAI21_X1 \mylsu/_1789_ ( .A(\mylsu/_0349_ ), .B1(\mylsu/_0383_ ), .B2(\mylsu/_0384_ ), .ZN(\mylsu/_0385_ ) );
OAI211_X2 \mylsu/_1790_ ( .A(\mylsu/_0385_ ), .B(\mylsu/_0354_ ), .C1(fanout_net_27 ), .C2(\mylsu/_0876_ ), .ZN(\mylsu/_0386_ ) );
OAI21_X1 \mylsu/_1791_ ( .A(\mylsu/_1016_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0387_ ) );
NAND2_X1 \mylsu/_1792_ ( .A1(\mylsu/_0386_ ), .A2(\mylsu/_0387_ ), .ZN(\mylsu/_0112_ ) );
INV_X4 \mylsu/_1793_ ( .A(\mylsu/_0349_ ), .ZN(\mylsu/_0388_ ) );
BUF_X8 \mylsu/_1794_ ( .A(\mylsu/_0388_ ), .Z(\mylsu/_0389_ ) );
MUX2_X1 \mylsu/_1795_ ( .A(\mylsu/_0830_ ), .B(\mylsu/_0812_ ), .S(\mylsu/_0693_ ), .Z(\mylsu/_0390_ ) );
NOR2_X1 \mylsu/_1796_ ( .A1(\mylsu/_0390_ ), .A2(\mylsu/_0706_ ), .ZN(\mylsu/_0391_ ) );
NOR3_X1 \mylsu/_1797_ ( .A1(\mylsu/_0687_ ), .A2(\mylsu/_0689_ ), .A3(\mylsu/_0812_ ), .ZN(\mylsu/_0392_ ) );
NOR3_X1 \mylsu/_1798_ ( .A1(\mylsu/_0391_ ), .A2(\mylsu/_0764_ ), .A3(\mylsu/_0392_ ), .ZN(\mylsu/_0393_ ) );
OAI221_X1 \mylsu/_1799_ ( .A(\mylsu/_0354_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0877_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0393_ ), .ZN(\mylsu/_0394_ ) );
OAI21_X1 \mylsu/_1800_ ( .A(\mylsu/_1017_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0395_ ) );
NAND2_X1 \mylsu/_1801_ ( .A1(\mylsu/_0394_ ), .A2(\mylsu/_0395_ ), .ZN(\mylsu/_0113_ ) );
INV_X1 \mylsu/_1802_ ( .A(\mylsu/_0687_ ), .ZN(\mylsu/_0396_ ) );
OAI21_X4 \mylsu/_1803_ ( .A(\mylsu/_0683_ ), .B1(\mylsu/_0390_ ), .B2(\mylsu/_0396_ ), .ZN(\mylsu/_0397_ ) );
BUF_X4 \mylsu/_1804_ ( .A(\mylsu/_0397_ ), .Z(\mylsu/_0398_ ) );
BUF_X4 \mylsu/_1805_ ( .A(\mylsu/_0689_ ), .Z(\mylsu/_0399_ ) );
BUF_X4 \mylsu/_1806_ ( .A(\mylsu/_0687_ ), .Z(\mylsu/_0400_ ) );
NOR2_X1 \mylsu/_1807_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0813_ ), .ZN(\mylsu/_0401_ ) );
NOR3_X1 \mylsu/_1808_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0401_ ), .ZN(\mylsu/_0402_ ) );
OAI221_X1 \mylsu/_1809_ ( .A(\mylsu/_0354_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0878_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0402_ ), .ZN(\mylsu/_0403_ ) );
OAI21_X1 \mylsu/_1810_ ( .A(\mylsu/_1018_ ), .B1(\mylsu/_0356_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0404_ ) );
NAND2_X1 \mylsu/_1811_ ( .A1(\mylsu/_0403_ ), .A2(\mylsu/_0404_ ), .ZN(\mylsu/_0114_ ) );
NOR2_X1 \mylsu/_1812_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0814_ ), .ZN(\mylsu/_0405_ ) );
NOR3_X1 \mylsu/_1813_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0405_ ), .ZN(\mylsu/_0406_ ) );
OAI221_X1 \mylsu/_1814_ ( .A(\mylsu/_0354_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0879_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0406_ ), .ZN(\mylsu/_0407_ ) );
BUF_X4 \mylsu/_1815_ ( .A(\mylsu/_0667_ ), .Z(\mylsu/_0408_ ) );
OAI21_X1 \mylsu/_1816_ ( .A(\mylsu/_1019_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0409_ ) );
NAND2_X1 \mylsu/_1817_ ( .A1(\mylsu/_0407_ ), .A2(\mylsu/_0409_ ), .ZN(\mylsu/_0115_ ) );
BUF_X4 \mylsu/_1818_ ( .A(\mylsu/_0699_ ), .Z(\mylsu/_0410_ ) );
NOR2_X1 \mylsu/_1819_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0815_ ), .ZN(\mylsu/_0411_ ) );
NOR3_X1 \mylsu/_1820_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0411_ ), .ZN(\mylsu/_0412_ ) );
OAI221_X1 \mylsu/_1821_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0880_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0412_ ), .ZN(\mylsu/_0413_ ) );
OAI21_X1 \mylsu/_1822_ ( .A(\mylsu/_1020_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0414_ ) );
NAND2_X1 \mylsu/_1823_ ( .A1(\mylsu/_0413_ ), .A2(\mylsu/_0414_ ), .ZN(\mylsu/_0116_ ) );
NOR2_X1 \mylsu/_1824_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0816_ ), .ZN(\mylsu/_0415_ ) );
NOR3_X1 \mylsu/_1825_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0415_ ), .ZN(\mylsu/_0416_ ) );
OAI221_X1 \mylsu/_1826_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0881_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0416_ ), .ZN(\mylsu/_0417_ ) );
OAI21_X1 \mylsu/_1827_ ( .A(\mylsu/_1021_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0418_ ) );
NAND2_X1 \mylsu/_1828_ ( .A1(\mylsu/_0417_ ), .A2(\mylsu/_0418_ ), .ZN(\mylsu/_0117_ ) );
NOR2_X1 \mylsu/_1829_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0818_ ), .ZN(\mylsu/_0419_ ) );
NOR3_X1 \mylsu/_1830_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0419_ ), .ZN(\mylsu/_0420_ ) );
OAI221_X1 \mylsu/_1831_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0883_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0420_ ), .ZN(\mylsu/_0421_ ) );
OAI21_X1 \mylsu/_1832_ ( .A(\mylsu/_1023_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0422_ ) );
NAND2_X1 \mylsu/_1833_ ( .A1(\mylsu/_0421_ ), .A2(\mylsu/_0422_ ), .ZN(\mylsu/_0118_ ) );
NOR2_X1 \mylsu/_1834_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0819_ ), .ZN(\mylsu/_0423_ ) );
NOR3_X1 \mylsu/_1835_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0423_ ), .ZN(\mylsu/_0424_ ) );
OAI221_X1 \mylsu/_1836_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0884_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0424_ ), .ZN(\mylsu/_0425_ ) );
OAI21_X1 \mylsu/_1837_ ( .A(\mylsu/_1024_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0426_ ) );
NAND2_X1 \mylsu/_1838_ ( .A1(\mylsu/_0425_ ), .A2(\mylsu/_0426_ ), .ZN(\mylsu/_0119_ ) );
NOR2_X1 \mylsu/_1839_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0820_ ), .ZN(\mylsu/_0427_ ) );
NOR3_X1 \mylsu/_1840_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0427_ ), .ZN(\mylsu/_0428_ ) );
OAI221_X1 \mylsu/_1841_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0885_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0428_ ), .ZN(\mylsu/_0429_ ) );
OAI21_X1 \mylsu/_1842_ ( .A(\mylsu/_1025_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0430_ ) );
NAND2_X1 \mylsu/_1843_ ( .A1(\mylsu/_0429_ ), .A2(\mylsu/_0430_ ), .ZN(\mylsu/_0120_ ) );
OR2_X4 \mylsu/_1844_ ( .A1(\mylsu/_0397_ ), .A2(\mylsu/_0689_ ), .ZN(\mylsu/_0431_ ) );
AOI21_X1 \mylsu/_1845_ ( .A(\mylsu/_0431_ ), .B1(\mylsu/_0767_ ), .B2(\mylsu/_0396_ ), .ZN(\mylsu/_0432_ ) );
OAI221_X1 \mylsu/_1846_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0886_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0432_ ), .ZN(\mylsu/_0433_ ) );
OAI21_X1 \mylsu/_1847_ ( .A(\mylsu/_1026_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0434_ ) );
NAND2_X1 \mylsu/_1848_ ( .A1(\mylsu/_0433_ ), .A2(\mylsu/_0434_ ), .ZN(\mylsu/_0121_ ) );
AOI21_X1 \mylsu/_1849_ ( .A(\mylsu/_0431_ ), .B1(\mylsu/_0675_ ), .B2(\mylsu/_0396_ ), .ZN(\mylsu/_0435_ ) );
OAI221_X1 \mylsu/_1850_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0887_ ), .C1(\mylsu/_0389_ ), .C2(\mylsu/_0435_ ), .ZN(\mylsu/_0436_ ) );
OAI21_X1 \mylsu/_1851_ ( .A(\mylsu/_1027_ ), .B1(\mylsu/_0408_ ), .B2(fanout_net_26 ), .ZN(\mylsu/_0437_ ) );
NAND2_X1 \mylsu/_1852_ ( .A1(\mylsu/_0436_ ), .A2(\mylsu/_0437_ ), .ZN(\mylsu/_0122_ ) );
NOR2_X1 \mylsu/_1853_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0823_ ), .ZN(\mylsu/_0438_ ) );
NOR3_X1 \mylsu/_1854_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0438_ ), .ZN(\mylsu/_0439_ ) );
OAI221_X1 \mylsu/_1855_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0888_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0439_ ), .ZN(\mylsu/_0440_ ) );
OAI21_X1 \mylsu/_1856_ ( .A(\mylsu/_1028_ ), .B1(\mylsu/_0408_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0441_ ) );
NAND2_X1 \mylsu/_1857_ ( .A1(\mylsu/_0440_ ), .A2(\mylsu/_0441_ ), .ZN(\mylsu/_0123_ ) );
NOR2_X1 \mylsu/_1858_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0824_ ), .ZN(\mylsu/_0442_ ) );
NOR3_X1 \mylsu/_1859_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0442_ ), .ZN(\mylsu/_0443_ ) );
OAI221_X1 \mylsu/_1860_ ( .A(\mylsu/_0410_ ), .B1(fanout_net_27 ), .B2(\mylsu/_0889_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0443_ ), .ZN(\mylsu/_0444_ ) );
OAI21_X1 \mylsu/_1861_ ( .A(\mylsu/_1029_ ), .B1(\mylsu/_0408_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0445_ ) );
NAND2_X1 \mylsu/_1862_ ( .A1(\mylsu/_0444_ ), .A2(\mylsu/_0445_ ), .ZN(\mylsu/_0124_ ) );
NOR2_X1 \mylsu/_1863_ ( .A1(\mylsu/_0400_ ), .A2(\mylsu/_0825_ ), .ZN(\mylsu/_0446_ ) );
NOR3_X1 \mylsu/_1864_ ( .A1(\mylsu/_0398_ ), .A2(\mylsu/_0399_ ), .A3(\mylsu/_0446_ ), .ZN(\mylsu/_0447_ ) );
OAI221_X1 \mylsu/_1865_ ( .A(\mylsu/_0410_ ), .B1(\mylsu/_0916_ ), .B2(\mylsu/_0890_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0447_ ), .ZN(\mylsu/_0448_ ) );
OAI21_X1 \mylsu/_1866_ ( .A(\mylsu/_1030_ ), .B1(\mylsu/_0668_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0449_ ) );
NAND2_X1 \mylsu/_1867_ ( .A1(\mylsu/_0448_ ), .A2(\mylsu/_0449_ ), .ZN(\mylsu/_0125_ ) );
NOR2_X1 \mylsu/_1868_ ( .A1(\mylsu/_0687_ ), .A2(\mylsu/_0826_ ), .ZN(\mylsu/_0450_ ) );
NOR3_X1 \mylsu/_1869_ ( .A1(\mylsu/_0397_ ), .A2(\mylsu/_0689_ ), .A3(\mylsu/_0450_ ), .ZN(\mylsu/_0451_ ) );
OAI221_X1 \mylsu/_1870_ ( .A(\mylsu/_0700_ ), .B1(\mylsu/_0916_ ), .B2(\mylsu/_0891_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0451_ ), .ZN(\mylsu/_0452_ ) );
OAI21_X1 \mylsu/_1871_ ( .A(\mylsu/_1031_ ), .B1(\mylsu/_0668_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0453_ ) );
NAND2_X1 \mylsu/_1872_ ( .A1(\mylsu/_0452_ ), .A2(\mylsu/_0453_ ), .ZN(\mylsu/_0126_ ) );
NOR2_X1 \mylsu/_1873_ ( .A1(\mylsu/_0687_ ), .A2(\mylsu/_0827_ ), .ZN(\mylsu/_0454_ ) );
NOR3_X1 \mylsu/_1874_ ( .A1(\mylsu/_0397_ ), .A2(\mylsu/_0689_ ), .A3(\mylsu/_0454_ ), .ZN(\mylsu/_0455_ ) );
OAI221_X1 \mylsu/_1875_ ( .A(\mylsu/_0700_ ), .B1(\mylsu/_0916_ ), .B2(\mylsu/_0892_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0455_ ), .ZN(\mylsu/_0456_ ) );
OAI21_X1 \mylsu/_1876_ ( .A(\mylsu/_1032_ ), .B1(\mylsu/_0668_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0457_ ) );
NAND2_X1 \mylsu/_1877_ ( .A1(\mylsu/_0456_ ), .A2(\mylsu/_0457_ ), .ZN(\mylsu/_0127_ ) );
NOR2_X1 \mylsu/_1878_ ( .A1(\mylsu/_0687_ ), .A2(\mylsu/_0829_ ), .ZN(\mylsu/_0458_ ) );
NOR3_X1 \mylsu/_1879_ ( .A1(\mylsu/_0397_ ), .A2(\mylsu/_0689_ ), .A3(\mylsu/_0458_ ), .ZN(\mylsu/_0459_ ) );
OAI221_X1 \mylsu/_1880_ ( .A(\mylsu/_0700_ ), .B1(\mylsu/_0916_ ), .B2(\mylsu/_0894_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0459_ ), .ZN(\mylsu/_0460_ ) );
OAI21_X1 \mylsu/_1881_ ( .A(\mylsu/_1034_ ), .B1(\mylsu/_0668_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0461_ ) );
NAND2_X1 \mylsu/_1882_ ( .A1(\mylsu/_0460_ ), .A2(\mylsu/_0461_ ), .ZN(\mylsu/_0128_ ) );
AOI21_X1 \mylsu/_1883_ ( .A(\mylsu/_0431_ ), .B1(\mylsu/_0761_ ), .B2(\mylsu/_0396_ ), .ZN(\mylsu/_0462_ ) );
OAI221_X1 \mylsu/_1884_ ( .A(\mylsu/_0700_ ), .B1(\mylsu/_0916_ ), .B2(\mylsu/_0895_ ), .C1(\mylsu/_0388_ ), .C2(\mylsu/_0462_ ), .ZN(\mylsu/_0463_ ) );
OAI21_X1 \mylsu/_1885_ ( .A(\mylsu/_1035_ ), .B1(\mylsu/_0668_ ), .B2(\mylsu/_0911_ ), .ZN(\mylsu/_0464_ ) );
NAND2_X1 \mylsu/_1886_ ( .A1(\mylsu/_0463_ ), .A2(\mylsu/_0464_ ), .ZN(\mylsu/_0129_ ) );
MUX2_X1 \mylsu/_1887_ ( .A(\mylsu/_0772_ ), .B(\mylsu/_0839_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0465_ ) );
MUX2_X1 \mylsu/_1888_ ( .A(\mylsu/_0979_ ), .B(\mylsu/_0465_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0132_ ) );
NAND3_X1 \mylsu/_1889_ ( .A1(\mylsu/_0646_ ), .A2(\mylsu/_0588_ ), .A3(\mylsu/_0647_ ), .ZN(\mylsu/_0466_ ) );
OAI211_X2 \mylsu/_1890_ ( .A(\mylsu/_0651_ ), .B(\mylsu/_0466_ ), .C1(\mylsu/_0783_ ), .C2(\mylsu/_0642_ ), .ZN(\mylsu/_0467_ ) );
OAI21_X1 \mylsu/_1891_ ( .A(\mylsu/_0990_ ), .B1(\mylsu/_0636_ ), .B2(\mylsu/_0649_ ), .ZN(\mylsu/_0468_ ) );
NAND2_X1 \mylsu/_1892_ ( .A1(\mylsu/_0467_ ), .A2(\mylsu/_0468_ ), .ZN(\mylsu/_0133_ ) );
MUX2_X1 \mylsu/_1893_ ( .A(\mylsu/_0794_ ), .B(\mylsu/_0861_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0469_ ) );
MUX2_X1 \mylsu/_1894_ ( .A(\mylsu/_1001_ ), .B(\mylsu/_0469_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0134_ ) );
MUX2_X1 \mylsu/_1895_ ( .A(\mylsu/_0797_ ), .B(\mylsu/_0864_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0470_ ) );
MUX2_X1 \mylsu/_1896_ ( .A(\mylsu/_1004_ ), .B(\mylsu/_0470_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0135_ ) );
MUX2_X1 \mylsu/_1897_ ( .A(\mylsu/_0798_ ), .B(\mylsu/_0865_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0471_ ) );
MUX2_X1 \mylsu/_1898_ ( .A(\mylsu/_1005_ ), .B(\mylsu/_0471_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0136_ ) );
MUX2_X1 \mylsu/_1899_ ( .A(\mylsu/_0799_ ), .B(\mylsu/_0866_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0472_ ) );
MUX2_X1 \mylsu/_1900_ ( .A(\mylsu/_1006_ ), .B(\mylsu/_0472_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0137_ ) );
MUX2_X1 \mylsu/_1901_ ( .A(\mylsu/_0800_ ), .B(\mylsu/_0867_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0473_ ) );
MUX2_X1 \mylsu/_1902_ ( .A(\mylsu/_1007_ ), .B(\mylsu/_0473_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0138_ ) );
MUX2_X1 \mylsu/_1903_ ( .A(\mylsu/_0801_ ), .B(\mylsu/_0868_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0474_ ) );
MUX2_X1 \mylsu/_1904_ ( .A(\mylsu/_1008_ ), .B(\mylsu/_0474_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0139_ ) );
MUX2_X1 \mylsu/_1905_ ( .A(\mylsu/_0802_ ), .B(\mylsu/_0869_ ), .S(\mylsu/_0642_ ), .Z(\mylsu/_0475_ ) );
MUX2_X1 \mylsu/_1906_ ( .A(\mylsu/_1009_ ), .B(\mylsu/_0475_ ), .S(\mylsu/_0664_ ), .Z(\mylsu/_0140_ ) );
BUF_X8 \mylsu/_1907_ ( .A(\mylsu/_0641_ ), .Z(\mylsu/_0476_ ) );
MUX2_X1 \mylsu/_1908_ ( .A(\mylsu/_0803_ ), .B(\mylsu/_0870_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0477_ ) );
BUF_X4 \mylsu/_1909_ ( .A(\mylsu/_0650_ ), .Z(\mylsu/_0478_ ) );
MUX2_X1 \mylsu/_1910_ ( .A(\mylsu/_1010_ ), .B(\mylsu/_0477_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0141_ ) );
MUX2_X1 \mylsu/_1911_ ( .A(\mylsu/_0773_ ), .B(\mylsu/_0840_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0479_ ) );
MUX2_X1 \mylsu/_1912_ ( .A(\mylsu/_0980_ ), .B(\mylsu/_0479_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0142_ ) );
MUX2_X1 \mylsu/_1913_ ( .A(\mylsu/_0774_ ), .B(\mylsu/_0841_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0480_ ) );
MUX2_X1 \mylsu/_1914_ ( .A(\mylsu/_0981_ ), .B(\mylsu/_0480_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0143_ ) );
MUX2_X1 \mylsu/_1915_ ( .A(\mylsu/_0775_ ), .B(\mylsu/_0842_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0481_ ) );
MUX2_X1 \mylsu/_1916_ ( .A(\mylsu/_0982_ ), .B(\mylsu/_0481_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0144_ ) );
MUX2_X1 \mylsu/_1917_ ( .A(\mylsu/_0776_ ), .B(\mylsu/_0843_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0482_ ) );
MUX2_X1 \mylsu/_1918_ ( .A(\mylsu/_0983_ ), .B(\mylsu/_0482_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0145_ ) );
MUX2_X1 \mylsu/_1919_ ( .A(\mylsu/_0777_ ), .B(\mylsu/_0844_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0483_ ) );
MUX2_X1 \mylsu/_1920_ ( .A(\mylsu/_0984_ ), .B(\mylsu/_0483_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0146_ ) );
MUX2_X1 \mylsu/_1921_ ( .A(\mylsu/_0778_ ), .B(\mylsu/_0845_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0484_ ) );
MUX2_X1 \mylsu/_1922_ ( .A(\mylsu/_0985_ ), .B(\mylsu/_0484_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0147_ ) );
MUX2_X1 \mylsu/_1923_ ( .A(\mylsu/_0779_ ), .B(\mylsu/_0846_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0485_ ) );
MUX2_X1 \mylsu/_1924_ ( .A(\mylsu/_0986_ ), .B(\mylsu/_0485_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0148_ ) );
MUX2_X1 \mylsu/_1925_ ( .A(\mylsu/_0780_ ), .B(\mylsu/_0847_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0486_ ) );
MUX2_X1 \mylsu/_1926_ ( .A(\mylsu/_0987_ ), .B(\mylsu/_0486_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0149_ ) );
MUX2_X1 \mylsu/_1927_ ( .A(\mylsu/_0781_ ), .B(\mylsu/_0848_ ), .S(\mylsu/_0476_ ), .Z(\mylsu/_0487_ ) );
MUX2_X1 \mylsu/_1928_ ( .A(\mylsu/_0988_ ), .B(\mylsu/_0487_ ), .S(\mylsu/_0478_ ), .Z(\mylsu/_0150_ ) );
BUF_X8 \mylsu/_1929_ ( .A(\mylsu/_0641_ ), .Z(\mylsu/_0488_ ) );
MUX2_X1 \mylsu/_1930_ ( .A(\mylsu/_0782_ ), .B(\mylsu/_0849_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0489_ ) );
BUF_X4 \mylsu/_1931_ ( .A(\mylsu/_0650_ ), .Z(\mylsu/_0490_ ) );
MUX2_X1 \mylsu/_1932_ ( .A(\mylsu/_0989_ ), .B(\mylsu/_0489_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0151_ ) );
MUX2_X1 \mylsu/_1933_ ( .A(\mylsu/_0784_ ), .B(\mylsu/_0851_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0491_ ) );
MUX2_X1 \mylsu/_1934_ ( .A(\mylsu/_0991_ ), .B(\mylsu/_0491_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0152_ ) );
MUX2_X1 \mylsu/_1935_ ( .A(\mylsu/_0785_ ), .B(\mylsu/_0852_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0492_ ) );
MUX2_X1 \mylsu/_1936_ ( .A(\mylsu/_0992_ ), .B(\mylsu/_0492_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0153_ ) );
MUX2_X1 \mylsu/_1937_ ( .A(\mylsu/_0786_ ), .B(\mylsu/_0853_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0493_ ) );
MUX2_X1 \mylsu/_1938_ ( .A(\mylsu/_0993_ ), .B(\mylsu/_0493_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0154_ ) );
MUX2_X1 \mylsu/_1939_ ( .A(\mylsu/_0787_ ), .B(\mylsu/_0854_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0494_ ) );
MUX2_X1 \mylsu/_1940_ ( .A(\mylsu/_0994_ ), .B(\mylsu/_0494_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0155_ ) );
MUX2_X1 \mylsu/_1941_ ( .A(\mylsu/_0788_ ), .B(\mylsu/_0855_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0495_ ) );
MUX2_X1 \mylsu/_1942_ ( .A(\mylsu/_0995_ ), .B(\mylsu/_0495_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0156_ ) );
MUX2_X1 \mylsu/_1943_ ( .A(\mylsu/_0789_ ), .B(\mylsu/_0856_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0496_ ) );
MUX2_X1 \mylsu/_1944_ ( .A(\mylsu/_0996_ ), .B(\mylsu/_0496_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0157_ ) );
MUX2_X1 \mylsu/_1945_ ( .A(\mylsu/_0790_ ), .B(\mylsu/_0857_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0497_ ) );
MUX2_X1 \mylsu/_1946_ ( .A(\mylsu/_0997_ ), .B(\mylsu/_0497_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0158_ ) );
MUX2_X1 \mylsu/_1947_ ( .A(\mylsu/_0791_ ), .B(\mylsu/_0858_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0498_ ) );
MUX2_X1 \mylsu/_1948_ ( .A(\mylsu/_0998_ ), .B(\mylsu/_0498_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0159_ ) );
MUX2_X1 \mylsu/_1949_ ( .A(\mylsu/_0792_ ), .B(\mylsu/_0859_ ), .S(\mylsu/_0488_ ), .Z(\mylsu/_0499_ ) );
MUX2_X1 \mylsu/_1950_ ( .A(\mylsu/_0999_ ), .B(\mylsu/_0499_ ), .S(\mylsu/_0490_ ), .Z(\mylsu/_0160_ ) );
MUX2_X1 \mylsu/_1951_ ( .A(\mylsu/_0793_ ), .B(\mylsu/_0860_ ), .S(\mylsu/_0641_ ), .Z(\mylsu/_0500_ ) );
MUX2_X1 \mylsu/_1952_ ( .A(\mylsu/_1000_ ), .B(\mylsu/_0500_ ), .S(\mylsu/_0650_ ), .Z(\mylsu/_0161_ ) );
MUX2_X1 \mylsu/_1953_ ( .A(\mylsu/_0795_ ), .B(\mylsu/_0862_ ), .S(\mylsu/_0641_ ), .Z(\mylsu/_0501_ ) );
MUX2_X1 \mylsu/_1954_ ( .A(\mylsu/_1002_ ), .B(\mylsu/_0501_ ), .S(\mylsu/_0650_ ), .Z(\mylsu/_0162_ ) );
MUX2_X1 \mylsu/_1955_ ( .A(\mylsu/_0796_ ), .B(\mylsu/_0863_ ), .S(\mylsu/_0641_ ), .Z(\mylsu/_0502_ ) );
MUX2_X1 \mylsu/_1956_ ( .A(\mylsu/_1003_ ), .B(\mylsu/_0502_ ), .S(\mylsu/_0650_ ), .Z(\mylsu/_0163_ ) );
AOI21_X1 \mylsu/_1957_ ( .A(\mylsu/_0645_ ), .B1(\mylsu/_0670_ ), .B2(\mylsu/_0649_ ), .ZN(\mylsu/_0164_ ) );
MUX2_X1 \mylsu/_1958_ ( .A(\mylsu/_0057_ ), .B(\mylsu/_0321_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0165_ ) );
MUX2_X1 \mylsu/_1959_ ( .A(\mylsu/_0068_ ), .B(\mylsu/_0332_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0166_ ) );
MUX2_X1 \mylsu/_1960_ ( .A(\mylsu/_0071_ ), .B(\mylsu/_0335_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0167_ ) );
MUX2_X1 \mylsu/_1961_ ( .A(\mylsu/_0072_ ), .B(\mylsu/_0336_ ), .S(\mylsu/_0633_ ), .Z(\mylsu/_0168_ ) );
BUF_X4 \mylsu/_1962_ ( .A(\mylsu/_0567_ ), .Z(\mylsu/_0503_ ) );
MUX2_X1 \mylsu/_1963_ ( .A(\mylsu/_0073_ ), .B(\mylsu/_0337_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0169_ ) );
MUX2_X1 \mylsu/_1964_ ( .A(\mylsu/_0074_ ), .B(\mylsu/_0338_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0170_ ) );
MUX2_X1 \mylsu/_1965_ ( .A(\mylsu/_0075_ ), .B(\mylsu/_0339_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0171_ ) );
MUX2_X1 \mylsu/_1966_ ( .A(\mylsu/_0076_ ), .B(\mylsu/_0340_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0172_ ) );
MUX2_X1 \mylsu/_1967_ ( .A(\mylsu/_0077_ ), .B(\mylsu/_0341_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0173_ ) );
MUX2_X1 \mylsu/_1968_ ( .A(\mylsu/_0047_ ), .B(\mylsu/_0311_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0174_ ) );
MUX2_X1 \mylsu/_1969_ ( .A(\mylsu/_0048_ ), .B(\mylsu/_0312_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0175_ ) );
MUX2_X1 \mylsu/_1970_ ( .A(\mylsu/_0049_ ), .B(\mylsu/_0313_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0176_ ) );
MUX2_X1 \mylsu/_1971_ ( .A(\mylsu/_0050_ ), .B(\mylsu/_0314_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0177_ ) );
MUX2_X1 \mylsu/_1972_ ( .A(\mylsu/_0051_ ), .B(\mylsu/_0315_ ), .S(\mylsu/_0503_ ), .Z(\mylsu/_0178_ ) );
BUF_X4 \mylsu/_1973_ ( .A(\mylsu/_0567_ ), .Z(\mylsu/_0504_ ) );
MUX2_X1 \mylsu/_1974_ ( .A(\mylsu/_0052_ ), .B(\mylsu/_0316_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0179_ ) );
MUX2_X1 \mylsu/_1975_ ( .A(\mylsu/_0053_ ), .B(\mylsu/_0317_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0180_ ) );
MUX2_X1 \mylsu/_1976_ ( .A(\mylsu/_0054_ ), .B(\mylsu/_0318_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0181_ ) );
MUX2_X1 \mylsu/_1977_ ( .A(\mylsu/_0055_ ), .B(\mylsu/_0319_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0182_ ) );
MUX2_X1 \mylsu/_1978_ ( .A(\mylsu/_0056_ ), .B(\mylsu/_0320_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0183_ ) );
MUX2_X1 \mylsu/_1979_ ( .A(\mylsu/_0058_ ), .B(\mylsu/_0322_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0184_ ) );
MUX2_X1 \mylsu/_1980_ ( .A(\mylsu/_0059_ ), .B(\mylsu/_0323_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0185_ ) );
MUX2_X1 \mylsu/_1981_ ( .A(\mylsu/_0060_ ), .B(\mylsu/_0324_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0186_ ) );
MUX2_X1 \mylsu/_1982_ ( .A(\mylsu/_0061_ ), .B(\mylsu/_0325_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0187_ ) );
MUX2_X1 \mylsu/_1983_ ( .A(\mylsu/_0062_ ), .B(\mylsu/_0326_ ), .S(\mylsu/_0504_ ), .Z(\mylsu/_0188_ ) );
BUF_X4 \mylsu/_1984_ ( .A(\mylsu/_0567_ ), .Z(\mylsu/_0505_ ) );
MUX2_X1 \mylsu/_1985_ ( .A(\mylsu/_0063_ ), .B(\mylsu/_0327_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0189_ ) );
MUX2_X1 \mylsu/_1986_ ( .A(\mylsu/_0064_ ), .B(\mylsu/_0328_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0190_ ) );
MUX2_X1 \mylsu/_1987_ ( .A(\mylsu/_0065_ ), .B(\mylsu/_0329_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0191_ ) );
MUX2_X1 \mylsu/_1988_ ( .A(\mylsu/_0066_ ), .B(\mylsu/_0330_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0192_ ) );
MUX2_X1 \mylsu/_1989_ ( .A(\mylsu/_0067_ ), .B(\mylsu/_0331_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0193_ ) );
MUX2_X1 \mylsu/_1990_ ( .A(\mylsu/_0069_ ), .B(\mylsu/_0333_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0194_ ) );
MUX2_X1 \mylsu/_1991_ ( .A(\mylsu/_0070_ ), .B(\mylsu/_0334_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0195_ ) );
NAND3_X1 \mylsu/_1992_ ( .A1(\mylsu/_0567_ ), .A2(\mylsu/_0536_ ), .A3(\mylsu/_0535_ ), .ZN(\mylsu/_0506_ ) );
NOR2_X4 \mylsu/_1993_ ( .A1(\mylsu/_0506_ ), .A2(\mylsu/_0561_ ), .ZN(\mylsu/_0507_ ) );
BUF_X4 \mylsu/_1994_ ( .A(\mylsu/_0507_ ), .Z(\mylsu/_0508_ ) );
MUX2_X1 \mylsu/_1995_ ( .A(\mylsu/_0266_ ), .B(\mylsu/_0310_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0196_ ) );
MUX2_X1 \mylsu/_1996_ ( .A(\mylsu/_0277_ ), .B(\mylsu/_0321_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0197_ ) );
MUX2_X1 \mylsu/_1997_ ( .A(\mylsu/_0288_ ), .B(\mylsu/_0332_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0198_ ) );
MUX2_X1 \mylsu/_1998_ ( .A(\mylsu/_0291_ ), .B(\mylsu/_0335_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0199_ ) );
MUX2_X1 \mylsu/_1999_ ( .A(\mylsu/_0292_ ), .B(\mylsu/_0336_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0200_ ) );
MUX2_X1 \mylsu/_2000_ ( .A(\mylsu/_0293_ ), .B(\mylsu/_0337_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0201_ ) );
MUX2_X1 \mylsu/_2001_ ( .A(\mylsu/_0294_ ), .B(\mylsu/_0338_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0202_ ) );
MUX2_X1 \mylsu/_2002_ ( .A(\mylsu/_0295_ ), .B(\mylsu/_0339_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0203_ ) );
MUX2_X1 \mylsu/_2003_ ( .A(\mylsu/_0296_ ), .B(\mylsu/_0340_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0204_ ) );
MUX2_X1 \mylsu/_2004_ ( .A(\mylsu/_0297_ ), .B(\mylsu/_0341_ ), .S(\mylsu/_0508_ ), .Z(\mylsu/_0205_ ) );
BUF_X4 \mylsu/_2005_ ( .A(\mylsu/_0507_ ), .Z(\mylsu/_0509_ ) );
MUX2_X1 \mylsu/_2006_ ( .A(\mylsu/_0267_ ), .B(\mylsu/_0311_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0206_ ) );
MUX2_X1 \mylsu/_2007_ ( .A(\mylsu/_0268_ ), .B(\mylsu/_0312_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0207_ ) );
MUX2_X1 \mylsu/_2008_ ( .A(\mylsu/_0269_ ), .B(\mylsu/_0313_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0208_ ) );
MUX2_X1 \mylsu/_2009_ ( .A(\mylsu/_0270_ ), .B(\mylsu/_0314_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0209_ ) );
MUX2_X1 \mylsu/_2010_ ( .A(\mylsu/_0271_ ), .B(\mylsu/_0315_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0210_ ) );
MUX2_X1 \mylsu/_2011_ ( .A(\mylsu/_0272_ ), .B(\mylsu/_0316_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0211_ ) );
MUX2_X1 \mylsu/_2012_ ( .A(\mylsu/_0273_ ), .B(\mylsu/_0317_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0212_ ) );
MUX2_X1 \mylsu/_2013_ ( .A(\mylsu/_0274_ ), .B(\mylsu/_0318_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0213_ ) );
MUX2_X1 \mylsu/_2014_ ( .A(\mylsu/_0275_ ), .B(\mylsu/_0319_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0214_ ) );
MUX2_X1 \mylsu/_2015_ ( .A(\mylsu/_0276_ ), .B(\mylsu/_0320_ ), .S(\mylsu/_0509_ ), .Z(\mylsu/_0215_ ) );
BUF_X4 \mylsu/_2016_ ( .A(\mylsu/_0507_ ), .Z(\mylsu/_0510_ ) );
MUX2_X1 \mylsu/_2017_ ( .A(\mylsu/_0278_ ), .B(\mylsu/_0322_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0216_ ) );
MUX2_X1 \mylsu/_2018_ ( .A(\mylsu/_0279_ ), .B(\mylsu/_0323_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0217_ ) );
MUX2_X1 \mylsu/_2019_ ( .A(\mylsu/_0280_ ), .B(\mylsu/_0324_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0218_ ) );
MUX2_X1 \mylsu/_2020_ ( .A(\mylsu/_0281_ ), .B(\mylsu/_0325_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0219_ ) );
MUX2_X1 \mylsu/_2021_ ( .A(\mylsu/_0282_ ), .B(\mylsu/_0326_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0220_ ) );
MUX2_X1 \mylsu/_2022_ ( .A(\mylsu/_0283_ ), .B(\mylsu/_0327_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0221_ ) );
MUX2_X1 \mylsu/_2023_ ( .A(\mylsu/_0284_ ), .B(\mylsu/_0328_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0222_ ) );
MUX2_X1 \mylsu/_2024_ ( .A(\mylsu/_0285_ ), .B(\mylsu/_0329_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0223_ ) );
MUX2_X1 \mylsu/_2025_ ( .A(\mylsu/_0286_ ), .B(\mylsu/_0330_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0224_ ) );
MUX2_X1 \mylsu/_2026_ ( .A(\mylsu/_0287_ ), .B(\mylsu/_0331_ ), .S(\mylsu/_0510_ ), .Z(\mylsu/_0225_ ) );
MUX2_X1 \mylsu/_2027_ ( .A(\mylsu/_0289_ ), .B(\mylsu/_0333_ ), .S(\mylsu/_0507_ ), .Z(\mylsu/_0226_ ) );
MUX2_X1 \mylsu/_2028_ ( .A(\mylsu/_0290_ ), .B(\mylsu/_0334_ ), .S(\mylsu/_0507_ ), .Z(\mylsu/_0227_ ) );
MUX2_X1 \mylsu/_2029_ ( .A(\mylsu/_0926_ ), .B(\mylsu/_0918_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0228_ ) );
MUX2_X1 \mylsu/_2030_ ( .A(\mylsu/_0927_ ), .B(\mylsu/_0919_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0229_ ) );
MUX2_X1 \mylsu/_2031_ ( .A(\mylsu/_0928_ ), .B(\mylsu/_0920_ ), .S(\mylsu/_0505_ ), .Z(\mylsu/_0230_ ) );
MUX2_X1 \mylsu/_2032_ ( .A(\mylsu/_0804_ ), .B(\mylsu/_0794_ ), .S(\mylsu/_0549_ ), .Z(\mylsu/_0511_ ) );
AND2_X1 \mylsu/_2033_ ( .A1(\mylsu/_0511_ ), .A2(\mylsu/_0531_ ), .ZN(\mylsu/_0080_ ) );
NAND3_X1 \mylsu/_2034_ ( .A1(\mylsu/_0541_ ), .A2(\mylsu/_0547_ ), .A3(\mylsu/_0563_ ), .ZN(\mylsu/_0512_ ) );
OAI21_X1 \mylsu/_2035_ ( .A(\mylsu/_0512_ ), .B1(\mylsu/_0546_ ), .B2(\mylsu/_0575_ ), .ZN(\mylsu/_0513_ ) );
NOR2_X1 \mylsu/_2036_ ( .A1(\mylsu/_0513_ ), .A2(\mylsu/_0564_ ), .ZN(\mylsu/_0514_ ) );
OAI21_X1 \mylsu/_2037_ ( .A(\mylsu/_0531_ ), .B1(\mylsu/_0514_ ), .B2(\mylsu/_1046_ ), .ZN(\mylsu/_0515_ ) );
NOR2_X1 \mylsu/_2038_ ( .A1(\mylsu/_0916_ ), .A2(\mylsu/_0914_ ), .ZN(\mylsu/_0516_ ) );
AND2_X1 \mylsu/_2039_ ( .A1(\mylsu/_0516_ ), .A2(\mylsu/_0929_ ), .ZN(\mylsu/_0517_ ) );
OAI211_X2 \mylsu/_2040_ ( .A(\mylsu/_0517_ ), .B(\mylsu/_0646_ ), .C1(\mylsu/_0534_ ), .C2(\mylsu/_0925_ ), .ZN(\mylsu/_0518_ ) );
AND2_X1 \mylsu/_2041_ ( .A1(\mylsu/_0518_ ), .A2(\mylsu/_0575_ ), .ZN(\mylsu/_0519_ ) );
AOI21_X1 \mylsu/_2042_ ( .A(\mylsu/_0515_ ), .B1(\mylsu/_0514_ ), .B2(\mylsu/_0519_ ), .ZN(\mylsu/_0130_ ) );
NAND2_X1 \mylsu/_2043_ ( .A1(\mylsu/_0356_ ), .A2(\mylsu/_0805_ ), .ZN(\mylsu/_0520_ ) );
OAI211_X2 \mylsu/_2044_ ( .A(\mylsu/_0546_ ), .B(\mylsu/_0916_ ), .C1(\mylsu/_0541_ ), .C2(\mylsu/_0929_ ), .ZN(\mylsu/_0521_ ) );
AOI21_X1 \mylsu/_2045_ ( .A(\mylsu/_0911_ ), .B1(\mylsu/_0520_ ), .B2(\mylsu/_0521_ ), .ZN(\mylsu/_0131_ ) );
OAI21_X1 \mylsu/_2046_ ( .A(\mylsu/_0531_ ), .B1(\mylsu/_0514_ ), .B2(\mylsu/_1043_ ), .ZN(\mylsu/_0522_ ) );
AND4_X1 \mylsu/_2047_ ( .A1(\mylsu/_0929_ ), .A2(\mylsu/_0923_ ), .A3(\mylsu/_0924_ ), .A4(\mylsu/_0925_ ), .ZN(\mylsu/_0523_ ) );
AND2_X1 \mylsu/_2048_ ( .A1(\mylsu/_0523_ ), .A2(\mylsu/_0516_ ), .ZN(\mylsu/_0524_ ) );
NOR3_X1 \mylsu/_2049_ ( .A1(\mylsu/_0513_ ), .A2(\mylsu/_0564_ ), .A3(\mylsu/_0524_ ), .ZN(\mylsu/_0525_ ) );
NOR2_X1 \mylsu/_2050_ ( .A1(\mylsu/_0522_ ), .A2(\mylsu/_0525_ ), .ZN(\mylsu/_0231_ ) );
OAI21_X1 \mylsu/_2051_ ( .A(\mylsu/_0531_ ), .B1(\mylsu/_0514_ ), .B2(\mylsu/_1044_ ), .ZN(\mylsu/_0526_ ) );
NAND3_X1 \mylsu/_2052_ ( .A1(\mylsu/_0517_ ), .A2(\mylsu/_0551_ ), .A3(\mylsu/_0634_ ), .ZN(\mylsu/_0527_ ) );
AOI21_X1 \mylsu/_2053_ ( .A(\mylsu/_0526_ ), .B1(\mylsu/_0525_ ), .B2(\mylsu/_0527_ ), .ZN(\mylsu/_0232_ ) );
NOR2_X1 \mylsu/_2054_ ( .A1(\mylsu/_0514_ ), .A2(\mylsu/_1045_ ), .ZN(\mylsu/_0528_ ) );
NAND4_X1 \mylsu/_2055_ ( .A1(\mylsu/_0516_ ), .A2(\mylsu/_0929_ ), .A3(\mylsu/_0924_ ), .A4(\mylsu/_0925_ ), .ZN(\mylsu/_0529_ ) );
AND2_X1 \mylsu/_2056_ ( .A1(\mylsu/_0527_ ), .A2(\mylsu/_0529_ ), .ZN(\mylsu/_0530_ ) );
AOI211_X2 \mylsu/_2057_ ( .A(\mylsu/_0911_ ), .B(\mylsu/_0528_ ), .C1(\mylsu/_0514_ ), .C2(\mylsu/_0530_ ), .ZN(\mylsu/_0233_ ) );
DFF_X1 \mylsu/_2058_ ( .D(\mylsu/_1212_ ), .CK(clock ), .Q(LS_WB_pc ), .QN(\mylsu/_1205_ ) );
DFF_X1 \mylsu/_2059_ ( .D(\mylsu/_1213_ ), .CK(clock ), .Q(\LS_WB_waddr_reg [0] ), .QN(\mylsu/_1204_ ) );
DFF_X1 \mylsu/_2060_ ( .D(\mylsu/_1214_ ), .CK(clock ), .Q(\LS_WB_waddr_reg [1] ), .QN(\mylsu/_1203_ ) );
DFF_X1 \mylsu/_2061_ ( .D(\mylsu/_1215_ ), .CK(clock ), .Q(\LS_WB_waddr_reg [2] ), .QN(\mylsu/_1202_ ) );
DFF_X1 \mylsu/_2062_ ( .D(\mylsu/_1216_ ), .CK(clock ), .Q(\LS_WB_waddr_reg [3] ), .QN(\mylsu/_1201_ ) );
DFF_X1 \mylsu/_2063_ ( .D(\mylsu/_1217_ ), .CK(clock ), .Q(\LS_WB_waddr_reg [4] ), .QN(\mylsu/_1200_ ) );
DFF_X1 \mylsu/_2064_ ( .D(\mylsu/_1218_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [0] ), .QN(\mylsu/_1199_ ) );
DFF_X1 \mylsu/_2065_ ( .D(\mylsu/_1219_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [1] ), .QN(\mylsu/_1198_ ) );
DFF_X1 \mylsu/_2066_ ( .D(\mylsu/_1220_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [2] ), .QN(\mylsu/_1197_ ) );
DFF_X1 \mylsu/_2067_ ( .D(\mylsu/_1221_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [3] ), .QN(\mylsu/_1196_ ) );
DFF_X1 \mylsu/_2068_ ( .D(\mylsu/_1222_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [4] ), .QN(\mylsu/_1195_ ) );
DFF_X1 \mylsu/_2069_ ( .D(\mylsu/_1223_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [5] ), .QN(\mylsu/_1194_ ) );
DFF_X1 \mylsu/_2070_ ( .D(\mylsu/_1224_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [6] ), .QN(\mylsu/_1193_ ) );
DFF_X1 \mylsu/_2071_ ( .D(\mylsu/_1225_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [7] ), .QN(\mylsu/_1192_ ) );
DFF_X1 \mylsu/_2072_ ( .D(\mylsu/_1226_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [8] ), .QN(\mylsu/_1191_ ) );
DFF_X1 \mylsu/_2073_ ( .D(\mylsu/_1227_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [9] ), .QN(\mylsu/_1190_ ) );
DFF_X1 \mylsu/_2074_ ( .D(\mylsu/_1228_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [10] ), .QN(\mylsu/_1189_ ) );
DFF_X1 \mylsu/_2075_ ( .D(\mylsu/_1229_ ), .CK(clock ), .Q(\LS_WB_waddr_csreg [11] ), .QN(\mylsu/_1188_ ) );
DFF_X1 \mylsu/_2076_ ( .D(\mylsu/_1230_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [0] ), .QN(\mylsu/_1187_ ) );
DFF_X1 \mylsu/_2077_ ( .D(\mylsu/_1231_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [1] ), .QN(\mylsu/_1186_ ) );
DFF_X1 \mylsu/_2078_ ( .D(\mylsu/_1232_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [2] ), .QN(\mylsu/_1185_ ) );
DFF_X1 \mylsu/_2079_ ( .D(\mylsu/_1233_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [3] ), .QN(\mylsu/_1184_ ) );
DFF_X1 \mylsu/_2080_ ( .D(\mylsu/_1234_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [4] ), .QN(\mylsu/_1183_ ) );
DFF_X1 \mylsu/_2081_ ( .D(\mylsu/_1235_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [5] ), .QN(\mylsu/_1182_ ) );
DFF_X1 \mylsu/_2082_ ( .D(\mylsu/_1236_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [6] ), .QN(\mylsu/_1181_ ) );
DFF_X1 \mylsu/_2083_ ( .D(\mylsu/_1237_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [7] ), .QN(\mylsu/_1180_ ) );
DFF_X1 \mylsu/_2084_ ( .D(\mylsu/_1238_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [8] ), .QN(\mylsu/_1179_ ) );
DFF_X1 \mylsu/_2085_ ( .D(\mylsu/_1239_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [9] ), .QN(\mylsu/_1178_ ) );
DFF_X1 \mylsu/_2086_ ( .D(\mylsu/_1240_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [10] ), .QN(\mylsu/_1177_ ) );
DFF_X1 \mylsu/_2087_ ( .D(\mylsu/_1241_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [11] ), .QN(\mylsu/_1176_ ) );
DFF_X1 \mylsu/_2088_ ( .D(\mylsu/_1242_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [12] ), .QN(\mylsu/_1175_ ) );
DFF_X1 \mylsu/_2089_ ( .D(\mylsu/_1243_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [13] ), .QN(\mylsu/_1174_ ) );
DFF_X1 \mylsu/_2090_ ( .D(\mylsu/_1244_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [14] ), .QN(\mylsu/_1173_ ) );
DFF_X1 \mylsu/_2091_ ( .D(\mylsu/_1245_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [15] ), .QN(\mylsu/_1172_ ) );
DFF_X1 \mylsu/_2092_ ( .D(\mylsu/_1246_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [16] ), .QN(\mylsu/_1171_ ) );
DFF_X1 \mylsu/_2093_ ( .D(\mylsu/_1247_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [17] ), .QN(\mylsu/_1170_ ) );
DFF_X1 \mylsu/_2094_ ( .D(\mylsu/_1248_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [18] ), .QN(\mylsu/_1169_ ) );
DFF_X1 \mylsu/_2095_ ( .D(\mylsu/_1249_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [19] ), .QN(\mylsu/_1168_ ) );
DFF_X1 \mylsu/_2096_ ( .D(\mylsu/_1250_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [20] ), .QN(\mylsu/_1167_ ) );
DFF_X1 \mylsu/_2097_ ( .D(\mylsu/_1251_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [21] ), .QN(\mylsu/_1166_ ) );
DFF_X1 \mylsu/_2098_ ( .D(\mylsu/_1252_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [22] ), .QN(\mylsu/_1165_ ) );
DFF_X1 \mylsu/_2099_ ( .D(\mylsu/_1253_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [23] ), .QN(\mylsu/_1164_ ) );
DFF_X1 \mylsu/_2100_ ( .D(\mylsu/_1254_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [24] ), .QN(\mylsu/_1163_ ) );
DFF_X1 \mylsu/_2101_ ( .D(\mylsu/_1255_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [25] ), .QN(\mylsu/_1162_ ) );
DFF_X1 \mylsu/_2102_ ( .D(\mylsu/_1256_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [26] ), .QN(\mylsu/_1161_ ) );
DFF_X1 \mylsu/_2103_ ( .D(\mylsu/_1257_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [27] ), .QN(\mylsu/_1160_ ) );
DFF_X1 \mylsu/_2104_ ( .D(\mylsu/_1258_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [28] ), .QN(\mylsu/_1159_ ) );
DFF_X1 \mylsu/_2105_ ( .D(\mylsu/_1259_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [29] ), .QN(\mylsu/_1158_ ) );
DFF_X1 \mylsu/_2106_ ( .D(\mylsu/_1260_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [30] ), .QN(\mylsu/_1157_ ) );
DFF_X1 \mylsu/_2107_ ( .D(\mylsu/_1261_ ), .CK(clock ), .Q(\LS_WB_wdata_reg [31] ), .QN(\mylsu/_1156_ ) );
DFF_X1 \mylsu/_2108_ ( .D(\mylsu/_1262_ ), .CK(clock ), .Q(LS_WB_wen_reg ), .QN(\mylsu/_1155_ ) );
DFF_X1 \mylsu/_2109_ ( .D(\mylsu/_1263_ ), .CK(clock ), .Q(previous_load_done ), .QN(\mylsu/_1154_ ) );
DFF_X1 \mylsu/_2110_ ( .D(\mylsu/_1264_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [0] ), .QN(\mylsu/_1153_ ) );
DFF_X1 \mylsu/_2111_ ( .D(\mylsu/_1265_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [1] ), .QN(\mylsu/_1152_ ) );
DFF_X1 \mylsu/_2112_ ( .D(\mylsu/_1266_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [2] ), .QN(\mylsu/_1151_ ) );
DFF_X1 \mylsu/_2113_ ( .D(\mylsu/_1267_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [3] ), .QN(\mylsu/_1150_ ) );
DFF_X1 \mylsu/_2114_ ( .D(\mylsu/_1268_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [4] ), .QN(\mylsu/_1149_ ) );
DFF_X1 \mylsu/_2115_ ( .D(\mylsu/_1269_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [5] ), .QN(\mylsu/_1148_ ) );
DFF_X1 \mylsu/_2116_ ( .D(\mylsu/_1270_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [6] ), .QN(\mylsu/_1147_ ) );
DFF_X1 \mylsu/_2117_ ( .D(\mylsu/_1271_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [7] ), .QN(\mylsu/_1146_ ) );
DFF_X1 \mylsu/_2118_ ( .D(\mylsu/_1272_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [8] ), .QN(\mylsu/_1145_ ) );
DFF_X1 \mylsu/_2119_ ( .D(\mylsu/_1273_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [9] ), .QN(\mylsu/_1144_ ) );
DFF_X1 \mylsu/_2120_ ( .D(\mylsu/_1274_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [10] ), .QN(\mylsu/_1143_ ) );
DFF_X1 \mylsu/_2121_ ( .D(\mylsu/_1275_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [11] ), .QN(\mylsu/_1142_ ) );
DFF_X1 \mylsu/_2122_ ( .D(\mylsu/_1276_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [12] ), .QN(\mylsu/_1141_ ) );
DFF_X1 \mylsu/_2123_ ( .D(\mylsu/_1277_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [13] ), .QN(\mylsu/_1140_ ) );
DFF_X1 \mylsu/_2124_ ( .D(\mylsu/_1278_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [14] ), .QN(\mylsu/_1139_ ) );
DFF_X1 \mylsu/_2125_ ( .D(\mylsu/_1279_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [15] ), .QN(\mylsu/_1138_ ) );
DFF_X1 \mylsu/_2126_ ( .D(\mylsu/_1280_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [16] ), .QN(\mylsu/_1137_ ) );
DFF_X1 \mylsu/_2127_ ( .D(\mylsu/_1281_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [17] ), .QN(\mylsu/_1136_ ) );
DFF_X1 \mylsu/_2128_ ( .D(\mylsu/_1282_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [18] ), .QN(\mylsu/_1135_ ) );
DFF_X1 \mylsu/_2129_ ( .D(\mylsu/_1283_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [19] ), .QN(\mylsu/_1134_ ) );
DFF_X1 \mylsu/_2130_ ( .D(\mylsu/_1284_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [20] ), .QN(\mylsu/_1133_ ) );
DFF_X1 \mylsu/_2131_ ( .D(\mylsu/_1285_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [21] ), .QN(\mylsu/_1132_ ) );
DFF_X1 \mylsu/_2132_ ( .D(\mylsu/_1286_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [22] ), .QN(\mylsu/_1131_ ) );
DFF_X1 \mylsu/_2133_ ( .D(\mylsu/_1287_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [23] ), .QN(\mylsu/_1130_ ) );
DFF_X1 \mylsu/_2134_ ( .D(\mylsu/_1288_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [24] ), .QN(\mylsu/_1129_ ) );
DFF_X1 \mylsu/_2135_ ( .D(\mylsu/_1289_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [25] ), .QN(\mylsu/_1128_ ) );
DFF_X1 \mylsu/_2136_ ( .D(\mylsu/_1290_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [26] ), .QN(\mylsu/_1127_ ) );
DFF_X1 \mylsu/_2137_ ( .D(\mylsu/_1291_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [27] ), .QN(\mylsu/_1126_ ) );
DFF_X1 \mylsu/_2138_ ( .D(\mylsu/_1292_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [28] ), .QN(\mylsu/_1125_ ) );
DFF_X1 \mylsu/_2139_ ( .D(\mylsu/_1293_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [29] ), .QN(\mylsu/_1124_ ) );
DFF_X1 \mylsu/_2140_ ( .D(\mylsu/_1294_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [30] ), .QN(\mylsu/_1123_ ) );
DFF_X1 \mylsu/_2141_ ( .D(\mylsu/_1295_ ), .CK(clock ), .Q(\LS_WB_wdata_csreg [31] ), .QN(\mylsu/_1122_ ) );
DFF_X1 \mylsu/_2142_ ( .D(\mylsu/_1296_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [0] ), .QN(\mylsu/_1121_ ) );
DFF_X1 \mylsu/_2143_ ( .D(\mylsu/_1297_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [1] ), .QN(\mylsu/_1120_ ) );
DFF_X1 \mylsu/_2144_ ( .D(\mylsu/_1298_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [2] ), .QN(\mylsu/_1119_ ) );
DFF_X1 \mylsu/_2145_ ( .D(\mylsu/_1299_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [3] ), .QN(\mylsu/_1118_ ) );
DFF_X1 \mylsu/_2146_ ( .D(\mylsu/_1300_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [4] ), .QN(\mylsu/_1117_ ) );
DFF_X1 \mylsu/_2147_ ( .D(\mylsu/_1301_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [5] ), .QN(\mylsu/_1116_ ) );
DFF_X1 \mylsu/_2148_ ( .D(\mylsu/_1302_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [6] ), .QN(\mylsu/_1115_ ) );
DFF_X1 \mylsu/_2149_ ( .D(\mylsu/_1303_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [7] ), .QN(\mylsu/_1114_ ) );
DFF_X1 \mylsu/_2150_ ( .D(\mylsu/_1304_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [8] ), .QN(\mylsu/_1113_ ) );
DFF_X1 \mylsu/_2151_ ( .D(\mylsu/_1305_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [9] ), .QN(\mylsu/_1112_ ) );
DFF_X1 \mylsu/_2152_ ( .D(\mylsu/_1306_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [10] ), .QN(\mylsu/_1111_ ) );
DFF_X1 \mylsu/_2153_ ( .D(\mylsu/_1307_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [11] ), .QN(\mylsu/_1110_ ) );
DFF_X1 \mylsu/_2154_ ( .D(\mylsu/_1308_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [12] ), .QN(\mylsu/_1109_ ) );
DFF_X1 \mylsu/_2155_ ( .D(\mylsu/_1309_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [13] ), .QN(\mylsu/_1108_ ) );
DFF_X1 \mylsu/_2156_ ( .D(\mylsu/_1310_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [14] ), .QN(\mylsu/_1107_ ) );
DFF_X1 \mylsu/_2157_ ( .D(\mylsu/_1311_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [15] ), .QN(\mylsu/_1106_ ) );
DFF_X1 \mylsu/_2158_ ( .D(\mylsu/_1312_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [16] ), .QN(\mylsu/_1105_ ) );
DFF_X1 \mylsu/_2159_ ( .D(\mylsu/_1313_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [17] ), .QN(\mylsu/_1104_ ) );
DFF_X1 \mylsu/_2160_ ( .D(\mylsu/_1314_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [18] ), .QN(\mylsu/_1103_ ) );
DFF_X1 \mylsu/_2161_ ( .D(\mylsu/_1315_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [19] ), .QN(\mylsu/_1102_ ) );
DFF_X1 \mylsu/_2162_ ( .D(\mylsu/_1316_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [20] ), .QN(\mylsu/_1101_ ) );
DFF_X1 \mylsu/_2163_ ( .D(\mylsu/_1317_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [21] ), .QN(\mylsu/_1100_ ) );
DFF_X1 \mylsu/_2164_ ( .D(\mylsu/_1318_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [22] ), .QN(\mylsu/_1099_ ) );
DFF_X1 \mylsu/_2165_ ( .D(\mylsu/_1319_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [23] ), .QN(\mylsu/_1098_ ) );
DFF_X1 \mylsu/_2166_ ( .D(\mylsu/_1320_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [24] ), .QN(\mylsu/_1097_ ) );
DFF_X1 \mylsu/_2167_ ( .D(\mylsu/_1321_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [25] ), .QN(\mylsu/_1096_ ) );
DFF_X1 \mylsu/_2168_ ( .D(\mylsu/_1322_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [26] ), .QN(\mylsu/_1095_ ) );
DFF_X1 \mylsu/_2169_ ( .D(\mylsu/_1323_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [27] ), .QN(\mylsu/_1094_ ) );
DFF_X1 \mylsu/_2170_ ( .D(\mylsu/_1324_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [28] ), .QN(\mylsu/_1093_ ) );
DFF_X1 \mylsu/_2171_ ( .D(\mylsu/_1325_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [29] ), .QN(\mylsu/_1092_ ) );
DFF_X1 \mylsu/_2172_ ( .D(\mylsu/_1326_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [30] ), .QN(\mylsu/_1091_ ) );
DFF_X1 \mylsu/_2173_ ( .D(\mylsu/_1327_ ), .CK(clock ), .Q(\mylsu/araddr_tmp [31] ), .QN(\mylsu/_1090_ ) );
DFF_X1 \mylsu/_2174_ ( .D(\mylsu/_1328_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [0] ), .QN(\mylsu/_1089_ ) );
DFF_X1 \mylsu/_2175_ ( .D(\mylsu/_1329_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [1] ), .QN(\mylsu/_1088_ ) );
DFF_X1 \mylsu/_2176_ ( .D(\mylsu/_1330_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [2] ), .QN(\mylsu/_1087_ ) );
DFF_X1 \mylsu/_2177_ ( .D(\mylsu/_1331_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [3] ), .QN(\mylsu/_1086_ ) );
DFF_X1 \mylsu/_2178_ ( .D(\mylsu/_1332_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [4] ), .QN(\mylsu/_1085_ ) );
DFF_X1 \mylsu/_2179_ ( .D(\mylsu/_1333_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [5] ), .QN(\mylsu/_1084_ ) );
DFF_X1 \mylsu/_2180_ ( .D(\mylsu/_1334_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [6] ), .QN(\mylsu/_1083_ ) );
DFF_X1 \mylsu/_2181_ ( .D(\mylsu/_1335_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [7] ), .QN(\mylsu/_1082_ ) );
DFF_X1 \mylsu/_2182_ ( .D(\mylsu/_1336_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [8] ), .QN(\mylsu/_1081_ ) );
DFF_X1 \mylsu/_2183_ ( .D(\mylsu/_1337_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [9] ), .QN(\mylsu/_1080_ ) );
DFF_X1 \mylsu/_2184_ ( .D(\mylsu/_1338_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [10] ), .QN(\mylsu/_1079_ ) );
DFF_X1 \mylsu/_2185_ ( .D(\mylsu/_1339_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [11] ), .QN(\mylsu/_1078_ ) );
DFF_X1 \mylsu/_2186_ ( .D(\mylsu/_1340_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [12] ), .QN(\mylsu/_1077_ ) );
DFF_X1 \mylsu/_2187_ ( .D(\mylsu/_1341_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [13] ), .QN(\mylsu/_1076_ ) );
DFF_X1 \mylsu/_2188_ ( .D(\mylsu/_1342_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [14] ), .QN(\mylsu/_1075_ ) );
DFF_X1 \mylsu/_2189_ ( .D(\mylsu/_1343_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [15] ), .QN(\mylsu/_1074_ ) );
DFF_X1 \mylsu/_2190_ ( .D(\mylsu/_1344_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [16] ), .QN(\mylsu/_1073_ ) );
DFF_X1 \mylsu/_2191_ ( .D(\mylsu/_1345_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [17] ), .QN(\mylsu/_1072_ ) );
DFF_X1 \mylsu/_2192_ ( .D(\mylsu/_1346_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [18] ), .QN(\mylsu/_1071_ ) );
DFF_X1 \mylsu/_2193_ ( .D(\mylsu/_1347_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [19] ), .QN(\mylsu/_1070_ ) );
DFF_X1 \mylsu/_2194_ ( .D(\mylsu/_1348_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [20] ), .QN(\mylsu/_1069_ ) );
DFF_X1 \mylsu/_2195_ ( .D(\mylsu/_1349_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [21] ), .QN(\mylsu/_1068_ ) );
DFF_X1 \mylsu/_2196_ ( .D(\mylsu/_1350_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [22] ), .QN(\mylsu/_1067_ ) );
DFF_X1 \mylsu/_2197_ ( .D(\mylsu/_1351_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [23] ), .QN(\mylsu/_1066_ ) );
DFF_X1 \mylsu/_2198_ ( .D(\mylsu/_1352_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [24] ), .QN(\mylsu/_1065_ ) );
DFF_X1 \mylsu/_2199_ ( .D(\mylsu/_1353_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [25] ), .QN(\mylsu/_1064_ ) );
DFF_X1 \mylsu/_2200_ ( .D(\mylsu/_1354_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [26] ), .QN(\mylsu/_1063_ ) );
DFF_X1 \mylsu/_2201_ ( .D(\mylsu/_1355_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [27] ), .QN(\mylsu/_1062_ ) );
DFF_X1 \mylsu/_2202_ ( .D(\mylsu/_1356_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [28] ), .QN(\mylsu/_1061_ ) );
DFF_X1 \mylsu/_2203_ ( .D(\mylsu/_1357_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [29] ), .QN(\mylsu/_1060_ ) );
DFF_X1 \mylsu/_2204_ ( .D(\mylsu/_1358_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [30] ), .QN(\mylsu/_1059_ ) );
DFF_X1 \mylsu/_2205_ ( .D(\mylsu/_1359_ ), .CK(clock ), .Q(\mylsu/awaddr_tmp [31] ), .QN(\mylsu/_1058_ ) );
DFF_X1 \mylsu/_2206_ ( .D(\mylsu/_1360_ ), .CK(clock ), .Q(\mylsu/typ_tmp [0] ), .QN(\mylsu/_1057_ ) );
DFF_X1 \mylsu/_2207_ ( .D(\mylsu/_1361_ ), .CK(clock ), .Q(\mylsu/typ_tmp [1] ), .QN(\mylsu/_1056_ ) );
DFF_X1 \mylsu/_2208_ ( .D(\mylsu/_1362_ ), .CK(clock ), .Q(\mylsu/typ_tmp [2] ), .QN(\mylsu/_0006_ ) );
DFF_X1 \mylsu/_2209_ ( .D(\mylsu/_1363_ ), .CK(clock ), .Q(\LS_WB_wen_csreg [3] ), .QN(\mylsu/_1055_ ) );
DFF_X1 \mylsu/_2210_ ( .D(\mylsu/_1364_ ), .CK(clock ), .Q(\LS_WB_wen_csreg [6] ), .QN(\mylsu/_1054_ ) );
DFF_X1 \mylsu/_2211_ ( .D(\mylsu/_1365_ ), .CK(clock ), .Q(\LS_WB_wen_csreg [7] ), .QN(\mylsu/_1206_ ) );
DFF_X1 \mylsu/_2212_ ( .D(\mylsu/_0000_ ), .CK(clock ), .Q(\mylsu/state [0] ), .QN(\mylsu/_0005_ ) );
DFF_X1 \mylsu/_2213_ ( .D(\mylsu/_0001_ ), .CK(clock ), .Q(\mylsu/state [1] ), .QN(\mylsu/_1207_ ) );
DFF_X1 \mylsu/_2214_ ( .D(\mylsu/_0002_ ), .CK(clock ), .Q(\mylsu/state [2] ), .QN(\mylsu/_1208_ ) );
DFF_X1 \mylsu/_2215_ ( .D(\mylsu/_0003_ ), .CK(clock ), .Q(\mylsu/state [3] ), .QN(\mylsu/_1209_ ) );
DFF_X1 \mylsu/_2216_ ( .D(\mylsu/_0004_ ), .CK(clock ), .Q(\mylsu/state [4] ), .QN(\mylsu/_1053_ ) );
LOGIC1_X1 \mylsu/_2217_ ( .Z(\mylsu/_1210_ ) );
LOGIC0_X1 \mylsu/_2218_ ( .Z(\mylsu/_1211_ ) );
BUF_X1 \mylsu/_2219_ ( .A(arready_LSU ), .Z(LSU_arready_set ) );
BUF_X1 \mylsu/_2220_ ( .A(awready_LSU ), .Z(LSU_awready_set ) );
BUF_X1 \mylsu/_2221_ ( .A(\mylsu/_1211_ ), .Z(\arburst_LSU [0] ) );
BUF_X1 \mylsu/_2222_ ( .A(\mylsu/_1211_ ), .Z(\arburst_LSU [1] ) );
BUF_X1 \mylsu/_2223_ ( .A(\mylsu/_1211_ ), .Z(\arid_LSU [0] ) );
BUF_X1 \mylsu/_2224_ ( .A(\mylsu/_1210_ ), .Z(\arid_LSU [1] ) );
BUF_X1 \mylsu/_2225_ ( .A(\mylsu/_1211_ ), .Z(\arid_LSU [2] ) );
BUF_X1 \mylsu/_2226_ ( .A(\mylsu/_1211_ ), .Z(\arid_LSU [3] ) );
BUF_X1 \mylsu/_2227_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [0] ) );
BUF_X1 \mylsu/_2228_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [1] ) );
BUF_X1 \mylsu/_2229_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [2] ) );
BUF_X1 \mylsu/_2230_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [3] ) );
BUF_X1 \mylsu/_2231_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [4] ) );
BUF_X1 \mylsu/_2232_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [5] ) );
BUF_X1 \mylsu/_2233_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [6] ) );
BUF_X1 \mylsu/_2234_ ( .A(\mylsu/_1211_ ), .Z(\arlen_LSU [7] ) );
BUF_X1 \mylsu/_2235_ ( .A(\EX_LS_typ [1] ), .Z(\arsize_LSU [0] ) );
BUF_X1 \mylsu/_2236_ ( .A(\EX_LS_typ [2] ), .Z(\arsize_LSU [1] ) );
BUF_X1 \mylsu/_2237_ ( .A(\EX_LS_typ [3] ), .Z(\arsize_LSU [2] ) );
BUF_X1 \mylsu/_2238_ ( .A(\mylsu/_1211_ ), .Z(\awburst_LSU [0] ) );
BUF_X1 \mylsu/_2239_ ( .A(\mylsu/_1211_ ), .Z(\awburst_LSU [1] ) );
BUF_X1 \mylsu/_2240_ ( .A(\mylsu/_1210_ ), .Z(\awid_LSU [0] ) );
BUF_X1 \mylsu/_2241_ ( .A(\mylsu/_1210_ ), .Z(\awid_LSU [1] ) );
BUF_X1 \mylsu/_2242_ ( .A(\mylsu/_1211_ ), .Z(\awid_LSU [2] ) );
BUF_X1 \mylsu/_2243_ ( .A(\mylsu/_1211_ ), .Z(\awid_LSU [3] ) );
BUF_X1 \mylsu/_2244_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [0] ) );
BUF_X1 \mylsu/_2245_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [1] ) );
BUF_X1 \mylsu/_2246_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [2] ) );
BUF_X1 \mylsu/_2247_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [3] ) );
BUF_X1 \mylsu/_2248_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [4] ) );
BUF_X1 \mylsu/_2249_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [5] ) );
BUF_X1 \mylsu/_2250_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [6] ) );
BUF_X1 \mylsu/_2251_ ( .A(\mylsu/_1211_ ), .Z(\awlen_LSU [7] ) );
BUF_X1 \mylsu/_2252_ ( .A(\mylsu/_1211_ ), .Z(\awsize_LSU [2] ) );
BUF_X1 \mylsu/_2253_ ( .A(rmem_quest_LSU ), .Z(rready_LSU ) );
BUF_X1 \mylsu/_2254_ ( .A(\LS_WB_wen_csreg [3] ), .Z(\LS_WB_wen_csreg [0] ) );
BUF_X1 \mylsu/_2255_ ( .A(\LS_WB_wen_csreg [6] ), .Z(\LS_WB_wen_csreg [1] ) );
BUF_X1 \mylsu/_2256_ ( .A(\mylsu/_1211_ ), .Z(\LS_WB_wen_csreg [2] ) );
BUF_X1 \mylsu/_2257_ ( .A(\mylsu/_1211_ ), .Z(\LS_WB_wen_csreg [4] ) );
BUF_X1 \mylsu/_2258_ ( .A(\mylsu/_1211_ ), .Z(\LS_WB_wen_csreg [5] ) );
BUF_X1 \mylsu/_2259_ ( .A(\mylsu/_1210_ ), .Z(wlast_LSU ) );
BUF_X1 \mylsu/_2260_ ( .A(\mylsu/state [0] ), .Z(\mylsu/_0913_ ) );
BUF_X1 \mylsu/_2261_ ( .A(EXU_valid_LSU ), .Z(\mylsu/_0929_ ) );
BUF_X1 \mylsu/_2262_ ( .A(reset ), .Z(\mylsu/_0911_ ) );
BUF_X1 \mylsu/_2263_ ( .A(\EX_LS_typ [5] ), .Z(\mylsu/_0923_ ) );
BUF_X1 \mylsu/_2264_ ( .A(\EX_LS_typ [6] ), .Z(\mylsu/_0924_ ) );
BUF_X1 \mylsu/_2265_ ( .A(\EX_LS_typ [7] ), .Z(\mylsu/_0925_ ) );
BUF_X1 \mylsu/_2266_ ( .A(wready_LSU ), .Z(\mylsu/_1047_ ) );
BUF_X1 \mylsu/_2267_ ( .A(awready_LSU ), .Z(\mylsu/_0298_ ) );
BUF_X1 \mylsu/_2268_ ( .A(\mylsu/state [3] ), .Z(\mylsu/_0916_ ) );
BUF_X1 \mylsu/_2269_ ( .A(\rresp_LSU [1] ), .Z(\mylsu/_0910_ ) );
BUF_X1 \mylsu/_2270_ ( .A(\rresp_LSU [0] ), .Z(\mylsu/_0909_ ) );
BUF_X1 \mylsu/_2271_ ( .A(rvalid_LSU ), .Z(\mylsu/_0912_ ) );
BUF_X1 \mylsu/_2272_ ( .A(rlast_LSU ), .Z(\mylsu/_0907_ ) );
BUF_X1 \mylsu/_2273_ ( .A(\rid_LSU [0] ), .Z(\mylsu/_0903_ ) );
BUF_X1 \mylsu/_2274_ ( .A(\rid_LSU [1] ), .Z(\mylsu/_0904_ ) );
BUF_X1 \mylsu/_2275_ ( .A(\rid_LSU [3] ), .Z(\mylsu/_0906_ ) );
BUF_X1 \mylsu/_2276_ ( .A(\rid_LSU [2] ), .Z(\mylsu/_0905_ ) );
BUF_X1 \mylsu/_2277_ ( .A(\mylsu/state [1] ), .Z(\mylsu/_0914_ ) );
BUF_X1 \mylsu/_2278_ ( .A(\bresp_LSU [1] ), .Z(\mylsu/_0308_ ) );
BUF_X1 \mylsu/_2279_ ( .A(\bresp_LSU [0] ), .Z(\mylsu/_0307_ ) );
BUF_X1 \mylsu/_2280_ ( .A(bvalid_LSU ), .Z(\mylsu/_0309_ ) );
BUF_X1 \mylsu/_2281_ ( .A(\bid_LSU [1] ), .Z(\mylsu/_0303_ ) );
BUF_X1 \mylsu/_2282_ ( .A(\bid_LSU [0] ), .Z(\mylsu/_0302_ ) );
BUF_X1 \mylsu/_2283_ ( .A(\bid_LSU [3] ), .Z(\mylsu/_0305_ ) );
BUF_X1 \mylsu/_2284_ ( .A(\bid_LSU [2] ), .Z(\mylsu/_0304_ ) );
BUF_X1 \mylsu/_2285_ ( .A(\mylsu/state [4] ), .Z(\mylsu/_0917_ ) );
BUF_X1 \mylsu/_2286_ ( .A(\mylsu/_0011_ ), .Z(\mylsu/_0004_ ) );
BUF_X1 \mylsu/_2287_ ( .A(arready_LSU ), .Z(\mylsu/_0078_ ) );
BUF_X1 \mylsu/_2288_ ( .A(\mylsu/_0010_ ), .Z(\mylsu/_0003_ ) );
BUF_X1 \mylsu/_2289_ ( .A(\mylsu/_0007_ ), .Z(\mylsu/_0000_ ) );
BUF_X1 \mylsu/_2290_ ( .A(\mylsu/state [2] ), .Z(\mylsu/_0915_ ) );
BUF_X1 \mylsu/_2291_ ( .A(\mylsu/_0008_ ), .Z(\mylsu/_0001_ ) );
BUF_X1 \mylsu/_2292_ ( .A(\mylsu/_0009_ ), .Z(\mylsu/_0002_ ) );
BUF_X1 \mylsu/_2293_ ( .A(\mylsu/_0005_ ), .Z(\mylsu/_0012_ ) );
BUF_X1 \mylsu/_2294_ ( .A(\mylsu/_0079_ ), .Z(arvalid_LSU ) );
BUF_X1 \mylsu/_2295_ ( .A(\mylsu/_0908_ ), .Z(rmem_quest_LSU ) );
BUF_X1 \mylsu/_2296_ ( .A(\mylsu/_0301_ ), .Z(awvalid_LSU ) );
BUF_X1 \mylsu/_2297_ ( .A(\mylsu/_1052_ ), .Z(wvalid_LSU ) );
BUF_X1 \mylsu/_2298_ ( .A(\mylsu/_0306_ ), .Z(bready_LSU ) );
BUF_X1 \mylsu/_2299_ ( .A(\mylsu/_0838_ ), .Z(LSU_ready_EXU ) );
BUF_X1 \mylsu/_2300_ ( .A(\EX_LS_result_csreg_mem [0] ), .Z(\mylsu/_0839_ ) );
BUF_X1 \mylsu/_2301_ ( .A(\EX_LS_pc [0] ), .Z(\mylsu/_0772_ ) );
BUF_X1 \mylsu/_2302_ ( .A(\EX_LS_result_csreg_mem [1] ), .Z(\mylsu/_0850_ ) );
BUF_X1 \mylsu/_2303_ ( .A(\EX_LS_pc [1] ), .Z(\mylsu/_0783_ ) );
BUF_X1 \mylsu/_2304_ ( .A(\EX_LS_result_csreg_mem [2] ), .Z(\mylsu/_0861_ ) );
BUF_X1 \mylsu/_2305_ ( .A(\EX_LS_pc [2] ), .Z(\mylsu/_0794_ ) );
BUF_X1 \mylsu/_2306_ ( .A(\EX_LS_result_csreg_mem [3] ), .Z(\mylsu/_0864_ ) );
BUF_X1 \mylsu/_2307_ ( .A(\EX_LS_pc [3] ), .Z(\mylsu/_0797_ ) );
BUF_X1 \mylsu/_2308_ ( .A(\EX_LS_result_csreg_mem [4] ), .Z(\mylsu/_0865_ ) );
BUF_X1 \mylsu/_2309_ ( .A(\EX_LS_pc [4] ), .Z(\mylsu/_0798_ ) );
BUF_X1 \mylsu/_2310_ ( .A(\EX_LS_result_csreg_mem [5] ), .Z(\mylsu/_0866_ ) );
BUF_X1 \mylsu/_2311_ ( .A(\EX_LS_pc [5] ), .Z(\mylsu/_0799_ ) );
BUF_X1 \mylsu/_2312_ ( .A(\EX_LS_result_csreg_mem [6] ), .Z(\mylsu/_0867_ ) );
BUF_X1 \mylsu/_2313_ ( .A(\EX_LS_pc [6] ), .Z(\mylsu/_0800_ ) );
BUF_X1 \mylsu/_2314_ ( .A(\EX_LS_result_csreg_mem [7] ), .Z(\mylsu/_0868_ ) );
BUF_X1 \mylsu/_2315_ ( .A(\EX_LS_pc [7] ), .Z(\mylsu/_0801_ ) );
BUF_X1 \mylsu/_2316_ ( .A(\EX_LS_result_csreg_mem [8] ), .Z(\mylsu/_0869_ ) );
BUF_X1 \mylsu/_2317_ ( .A(\EX_LS_pc [8] ), .Z(\mylsu/_0802_ ) );
BUF_X1 \mylsu/_2318_ ( .A(\EX_LS_result_csreg_mem [9] ), .Z(\mylsu/_0870_ ) );
BUF_X1 \mylsu/_2319_ ( .A(\EX_LS_pc [9] ), .Z(\mylsu/_0803_ ) );
BUF_X1 \mylsu/_2320_ ( .A(\EX_LS_result_csreg_mem [10] ), .Z(\mylsu/_0840_ ) );
BUF_X1 \mylsu/_2321_ ( .A(\EX_LS_pc [10] ), .Z(\mylsu/_0773_ ) );
BUF_X1 \mylsu/_2322_ ( .A(\EX_LS_result_csreg_mem [11] ), .Z(\mylsu/_0841_ ) );
BUF_X1 \mylsu/_2323_ ( .A(\EX_LS_pc [11] ), .Z(\mylsu/_0774_ ) );
BUF_X1 \mylsu/_2324_ ( .A(\EX_LS_result_csreg_mem [12] ), .Z(\mylsu/_0842_ ) );
BUF_X1 \mylsu/_2325_ ( .A(\EX_LS_pc [12] ), .Z(\mylsu/_0775_ ) );
BUF_X1 \mylsu/_2326_ ( .A(\EX_LS_result_csreg_mem [13] ), .Z(\mylsu/_0843_ ) );
BUF_X1 \mylsu/_2327_ ( .A(\EX_LS_pc [13] ), .Z(\mylsu/_0776_ ) );
BUF_X1 \mylsu/_2328_ ( .A(\EX_LS_result_csreg_mem [14] ), .Z(\mylsu/_0844_ ) );
BUF_X1 \mylsu/_2329_ ( .A(\EX_LS_pc [14] ), .Z(\mylsu/_0777_ ) );
BUF_X1 \mylsu/_2330_ ( .A(\EX_LS_result_csreg_mem [15] ), .Z(\mylsu/_0845_ ) );
BUF_X1 \mylsu/_2331_ ( .A(\EX_LS_pc [15] ), .Z(\mylsu/_0778_ ) );
BUF_X1 \mylsu/_2332_ ( .A(\EX_LS_result_csreg_mem [16] ), .Z(\mylsu/_0846_ ) );
BUF_X1 \mylsu/_2333_ ( .A(\EX_LS_pc [16] ), .Z(\mylsu/_0779_ ) );
BUF_X1 \mylsu/_2334_ ( .A(\EX_LS_result_csreg_mem [17] ), .Z(\mylsu/_0847_ ) );
BUF_X1 \mylsu/_2335_ ( .A(\EX_LS_pc [17] ), .Z(\mylsu/_0780_ ) );
BUF_X1 \mylsu/_2336_ ( .A(\EX_LS_result_csreg_mem [18] ), .Z(\mylsu/_0848_ ) );
BUF_X1 \mylsu/_2337_ ( .A(\EX_LS_pc [18] ), .Z(\mylsu/_0781_ ) );
BUF_X1 \mylsu/_2338_ ( .A(\EX_LS_result_csreg_mem [19] ), .Z(\mylsu/_0849_ ) );
BUF_X1 \mylsu/_2339_ ( .A(\EX_LS_pc [19] ), .Z(\mylsu/_0782_ ) );
BUF_X1 \mylsu/_2340_ ( .A(\EX_LS_result_csreg_mem [20] ), .Z(\mylsu/_0851_ ) );
BUF_X1 \mylsu/_2341_ ( .A(\EX_LS_pc [20] ), .Z(\mylsu/_0784_ ) );
BUF_X1 \mylsu/_2342_ ( .A(\EX_LS_result_csreg_mem [21] ), .Z(\mylsu/_0852_ ) );
BUF_X1 \mylsu/_2343_ ( .A(\EX_LS_pc [21] ), .Z(\mylsu/_0785_ ) );
BUF_X1 \mylsu/_2344_ ( .A(\EX_LS_result_csreg_mem [22] ), .Z(\mylsu/_0853_ ) );
BUF_X1 \mylsu/_2345_ ( .A(\EX_LS_pc [22] ), .Z(\mylsu/_0786_ ) );
BUF_X1 \mylsu/_2346_ ( .A(\EX_LS_result_csreg_mem [23] ), .Z(\mylsu/_0854_ ) );
BUF_X1 \mylsu/_2347_ ( .A(\EX_LS_pc [23] ), .Z(\mylsu/_0787_ ) );
BUF_X1 \mylsu/_2348_ ( .A(\EX_LS_result_csreg_mem [24] ), .Z(\mylsu/_0855_ ) );
BUF_X1 \mylsu/_2349_ ( .A(\EX_LS_pc [24] ), .Z(\mylsu/_0788_ ) );
BUF_X1 \mylsu/_2350_ ( .A(\EX_LS_result_csreg_mem [25] ), .Z(\mylsu/_0856_ ) );
BUF_X1 \mylsu/_2351_ ( .A(\EX_LS_pc [25] ), .Z(\mylsu/_0789_ ) );
BUF_X1 \mylsu/_2352_ ( .A(\EX_LS_result_csreg_mem [26] ), .Z(\mylsu/_0857_ ) );
BUF_X1 \mylsu/_2353_ ( .A(\EX_LS_pc [26] ), .Z(\mylsu/_0790_ ) );
BUF_X1 \mylsu/_2354_ ( .A(\EX_LS_result_csreg_mem [27] ), .Z(\mylsu/_0858_ ) );
BUF_X1 \mylsu/_2355_ ( .A(\EX_LS_pc [27] ), .Z(\mylsu/_0791_ ) );
BUF_X1 \mylsu/_2356_ ( .A(\EX_LS_result_csreg_mem [28] ), .Z(\mylsu/_0859_ ) );
BUF_X1 \mylsu/_2357_ ( .A(\EX_LS_pc [28] ), .Z(\mylsu/_0792_ ) );
BUF_X1 \mylsu/_2358_ ( .A(\EX_LS_result_csreg_mem [29] ), .Z(\mylsu/_0860_ ) );
BUF_X1 \mylsu/_2359_ ( .A(\EX_LS_pc [29] ), .Z(\mylsu/_0793_ ) );
BUF_X1 \mylsu/_2360_ ( .A(\EX_LS_result_csreg_mem [30] ), .Z(\mylsu/_0862_ ) );
BUF_X1 \mylsu/_2361_ ( .A(\EX_LS_pc [30] ), .Z(\mylsu/_0795_ ) );
BUF_X1 \mylsu/_2362_ ( .A(\EX_LS_result_csreg_mem [31] ), .Z(\mylsu/_0863_ ) );
BUF_X1 \mylsu/_2363_ ( .A(\EX_LS_pc [31] ), .Z(\mylsu/_0796_ ) );
BUF_X1 \mylsu/_2364_ ( .A(\mylsu/araddr_tmp [0] ), .Z(\mylsu/_0046_ ) );
BUF_X1 \mylsu/_2365_ ( .A(\mylsu/araddr_tmp [1] ), .Z(\mylsu/_0057_ ) );
BUF_X1 \mylsu/_2366_ ( .A(\rdata_LSU [24] ), .Z(\mylsu/_0822_ ) );
BUF_X1 \mylsu/_2367_ ( .A(\rdata_LSU [16] ), .Z(\mylsu/_0813_ ) );
BUF_X1 \mylsu/_2368_ ( .A(\rdata_LSU [8] ), .Z(\mylsu/_0836_ ) );
BUF_X1 \mylsu/_2369_ ( .A(\rdata_LSU [0] ), .Z(\mylsu/_0806_ ) );
BUF_X1 \mylsu/_2370_ ( .A(\mylsu/typ_tmp [1] ), .Z(\mylsu/_0927_ ) );
BUF_X1 \mylsu/_2371_ ( .A(\mylsu/typ_tmp [0] ), .Z(\mylsu/_0926_ ) );
BUF_X1 \mylsu/_2372_ ( .A(\mylsu/_0006_ ), .Z(\mylsu/_0013_ ) );
BUF_X1 \mylsu/_2373_ ( .A(\mylsu/typ_tmp [2] ), .Z(\mylsu/_0928_ ) );
BUF_X1 \mylsu/_2374_ ( .A(\EX_LS_result_reg [0] ), .Z(\mylsu/_0871_ ) );
BUF_X1 \mylsu/_2375_ ( .A(\rdata_LSU [25] ), .Z(\mylsu/_0823_ ) );
BUF_X1 \mylsu/_2376_ ( .A(\rdata_LSU [17] ), .Z(\mylsu/_0814_ ) );
BUF_X1 \mylsu/_2377_ ( .A(\rdata_LSU [9] ), .Z(\mylsu/_0837_ ) );
BUF_X1 \mylsu/_2378_ ( .A(\rdata_LSU [1] ), .Z(\mylsu/_0817_ ) );
BUF_X1 \mylsu/_2379_ ( .A(\EX_LS_result_reg [1] ), .Z(\mylsu/_0882_ ) );
BUF_X1 \mylsu/_2380_ ( .A(\rdata_LSU [26] ), .Z(\mylsu/_0824_ ) );
BUF_X1 \mylsu/_2381_ ( .A(\rdata_LSU [18] ), .Z(\mylsu/_0815_ ) );
BUF_X1 \mylsu/_2382_ ( .A(\rdata_LSU [10] ), .Z(\mylsu/_0807_ ) );
BUF_X1 \mylsu/_2383_ ( .A(\rdata_LSU [2] ), .Z(\mylsu/_0828_ ) );
BUF_X1 \mylsu/_2384_ ( .A(\EX_LS_result_reg [2] ), .Z(\mylsu/_0893_ ) );
BUF_X1 \mylsu/_2385_ ( .A(\rdata_LSU [27] ), .Z(\mylsu/_0825_ ) );
BUF_X1 \mylsu/_2386_ ( .A(\rdata_LSU [19] ), .Z(\mylsu/_0816_ ) );
BUF_X1 \mylsu/_2387_ ( .A(\rdata_LSU [11] ), .Z(\mylsu/_0808_ ) );
BUF_X1 \mylsu/_2388_ ( .A(\rdata_LSU [3] ), .Z(\mylsu/_0831_ ) );
BUF_X1 \mylsu/_2389_ ( .A(\EX_LS_result_reg [3] ), .Z(\mylsu/_0896_ ) );
BUF_X1 \mylsu/_2390_ ( .A(\rdata_LSU [28] ), .Z(\mylsu/_0826_ ) );
BUF_X1 \mylsu/_2391_ ( .A(\rdata_LSU [20] ), .Z(\mylsu/_0818_ ) );
BUF_X1 \mylsu/_2392_ ( .A(\rdata_LSU [12] ), .Z(\mylsu/_0809_ ) );
BUF_X1 \mylsu/_2393_ ( .A(\rdata_LSU [4] ), .Z(\mylsu/_0832_ ) );
BUF_X1 \mylsu/_2394_ ( .A(\EX_LS_result_reg [4] ), .Z(\mylsu/_0897_ ) );
BUF_X1 \mylsu/_2395_ ( .A(\rdata_LSU [29] ), .Z(\mylsu/_0827_ ) );
BUF_X1 \mylsu/_2396_ ( .A(\rdata_LSU [21] ), .Z(\mylsu/_0819_ ) );
BUF_X1 \mylsu/_2397_ ( .A(\rdata_LSU [13] ), .Z(\mylsu/_0810_ ) );
BUF_X1 \mylsu/_2398_ ( .A(\rdata_LSU [5] ), .Z(\mylsu/_0833_ ) );
BUF_X1 \mylsu/_2399_ ( .A(\EX_LS_result_reg [5] ), .Z(\mylsu/_0898_ ) );
BUF_X1 \mylsu/_2400_ ( .A(\rdata_LSU [30] ), .Z(\mylsu/_0829_ ) );
BUF_X1 \mylsu/_2401_ ( .A(\rdata_LSU [22] ), .Z(\mylsu/_0820_ ) );
BUF_X1 \mylsu/_2402_ ( .A(\rdata_LSU [14] ), .Z(\mylsu/_0811_ ) );
BUF_X1 \mylsu/_2403_ ( .A(\rdata_LSU [6] ), .Z(\mylsu/_0834_ ) );
BUF_X1 \mylsu/_2404_ ( .A(\EX_LS_result_reg [6] ), .Z(\mylsu/_0899_ ) );
BUF_X1 \mylsu/_2405_ ( .A(\rdata_LSU [31] ), .Z(\mylsu/_0830_ ) );
BUF_X1 \mylsu/_2406_ ( .A(\rdata_LSU [23] ), .Z(\mylsu/_0821_ ) );
BUF_X1 \mylsu/_2407_ ( .A(\rdata_LSU [15] ), .Z(\mylsu/_0812_ ) );
BUF_X1 \mylsu/_2408_ ( .A(\rdata_LSU [7] ), .Z(\mylsu/_0835_ ) );
BUF_X1 \mylsu/_2409_ ( .A(\EX_LS_result_reg [7] ), .Z(\mylsu/_0900_ ) );
BUF_X1 \mylsu/_2410_ ( .A(\EX_LS_result_reg [8] ), .Z(\mylsu/_0901_ ) );
BUF_X1 \mylsu/_2411_ ( .A(\EX_LS_result_reg [9] ), .Z(\mylsu/_0902_ ) );
BUF_X1 \mylsu/_2412_ ( .A(\EX_LS_result_reg [10] ), .Z(\mylsu/_0872_ ) );
BUF_X1 \mylsu/_2413_ ( .A(\EX_LS_result_reg [11] ), .Z(\mylsu/_0873_ ) );
BUF_X1 \mylsu/_2414_ ( .A(\EX_LS_result_reg [12] ), .Z(\mylsu/_0874_ ) );
BUF_X1 \mylsu/_2415_ ( .A(\EX_LS_result_reg [13] ), .Z(\mylsu/_0875_ ) );
BUF_X1 \mylsu/_2416_ ( .A(\EX_LS_result_reg [14] ), .Z(\mylsu/_0876_ ) );
BUF_X1 \mylsu/_2417_ ( .A(\EX_LS_result_reg [15] ), .Z(\mylsu/_0877_ ) );
BUF_X1 \mylsu/_2418_ ( .A(\EX_LS_result_reg [16] ), .Z(\mylsu/_0878_ ) );
BUF_X1 \mylsu/_2419_ ( .A(\EX_LS_result_reg [17] ), .Z(\mylsu/_0879_ ) );
BUF_X1 \mylsu/_2420_ ( .A(\EX_LS_result_reg [18] ), .Z(\mylsu/_0880_ ) );
BUF_X1 \mylsu/_2421_ ( .A(\EX_LS_result_reg [19] ), .Z(\mylsu/_0881_ ) );
BUF_X1 \mylsu/_2422_ ( .A(\EX_LS_result_reg [20] ), .Z(\mylsu/_0883_ ) );
BUF_X1 \mylsu/_2423_ ( .A(\EX_LS_result_reg [21] ), .Z(\mylsu/_0884_ ) );
BUF_X1 \mylsu/_2424_ ( .A(\EX_LS_result_reg [22] ), .Z(\mylsu/_0885_ ) );
BUF_X1 \mylsu/_2425_ ( .A(\EX_LS_result_reg [23] ), .Z(\mylsu/_0886_ ) );
BUF_X1 \mylsu/_2426_ ( .A(\EX_LS_result_reg [24] ), .Z(\mylsu/_0887_ ) );
BUF_X1 \mylsu/_2427_ ( .A(\EX_LS_result_reg [25] ), .Z(\mylsu/_0888_ ) );
BUF_X1 \mylsu/_2428_ ( .A(\EX_LS_result_reg [26] ), .Z(\mylsu/_0889_ ) );
BUF_X1 \mylsu/_2429_ ( .A(\EX_LS_result_reg [27] ), .Z(\mylsu/_0890_ ) );
BUF_X1 \mylsu/_2430_ ( .A(\EX_LS_result_reg [28] ), .Z(\mylsu/_0891_ ) );
BUF_X1 \mylsu/_2431_ ( .A(\EX_LS_result_reg [29] ), .Z(\mylsu/_0892_ ) );
BUF_X1 \mylsu/_2432_ ( .A(\EX_LS_result_reg [30] ), .Z(\mylsu/_0894_ ) );
BUF_X1 \mylsu/_2433_ ( .A(\EX_LS_result_reg [31] ), .Z(\mylsu/_0895_ ) );
BUF_X1 \mylsu/_2434_ ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(\mylsu/_0310_ ) );
BUF_X1 \mylsu/_2435_ ( .A(\mylsu/_0014_ ), .Z(\araddr_LSU [0] ) );
BUF_X1 \mylsu/_2436_ ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(\mylsu/_0321_ ) );
BUF_X1 \mylsu/_2437_ ( .A(\mylsu/_0025_ ), .Z(\araddr_LSU [1] ) );
BUF_X1 \mylsu/_2438_ ( .A(\mylsu/araddr_tmp [2] ), .Z(\mylsu/_0068_ ) );
BUF_X1 \mylsu/_2439_ ( .A(\EX_LS_dest_csreg_mem [2] ), .Z(\mylsu/_0332_ ) );
BUF_X1 \mylsu/_2440_ ( .A(\mylsu/_0036_ ), .Z(\araddr_LSU [2] ) );
BUF_X1 \mylsu/_2441_ ( .A(\mylsu/araddr_tmp [3] ), .Z(\mylsu/_0071_ ) );
BUF_X1 \mylsu/_2442_ ( .A(\EX_LS_dest_csreg_mem [3] ), .Z(\mylsu/_0335_ ) );
BUF_X1 \mylsu/_2443_ ( .A(\mylsu/_0039_ ), .Z(\araddr_LSU [3] ) );
BUF_X1 \mylsu/_2444_ ( .A(\mylsu/araddr_tmp [4] ), .Z(\mylsu/_0072_ ) );
BUF_X1 \mylsu/_2445_ ( .A(\EX_LS_dest_csreg_mem [4] ), .Z(\mylsu/_0336_ ) );
BUF_X1 \mylsu/_2446_ ( .A(\mylsu/_0040_ ), .Z(\araddr_LSU [4] ) );
BUF_X1 \mylsu/_2447_ ( .A(\mylsu/araddr_tmp [5] ), .Z(\mylsu/_0073_ ) );
BUF_X1 \mylsu/_2448_ ( .A(\EX_LS_dest_csreg_mem [5] ), .Z(\mylsu/_0337_ ) );
BUF_X1 \mylsu/_2449_ ( .A(\mylsu/_0041_ ), .Z(\araddr_LSU [5] ) );
BUF_X1 \mylsu/_2450_ ( .A(\mylsu/araddr_tmp [6] ), .Z(\mylsu/_0074_ ) );
BUF_X1 \mylsu/_2451_ ( .A(\EX_LS_dest_csreg_mem [6] ), .Z(\mylsu/_0338_ ) );
BUF_X1 \mylsu/_2452_ ( .A(\mylsu/_0042_ ), .Z(\araddr_LSU [6] ) );
BUF_X1 \mylsu/_2453_ ( .A(\mylsu/araddr_tmp [7] ), .Z(\mylsu/_0075_ ) );
BUF_X1 \mylsu/_2454_ ( .A(\EX_LS_dest_csreg_mem [7] ), .Z(\mylsu/_0339_ ) );
BUF_X1 \mylsu/_2455_ ( .A(\mylsu/_0043_ ), .Z(\araddr_LSU [7] ) );
BUF_X1 \mylsu/_2456_ ( .A(\mylsu/araddr_tmp [8] ), .Z(\mylsu/_0076_ ) );
BUF_X1 \mylsu/_2457_ ( .A(\EX_LS_dest_csreg_mem [8] ), .Z(\mylsu/_0340_ ) );
BUF_X1 \mylsu/_2458_ ( .A(\mylsu/_0044_ ), .Z(\araddr_LSU [8] ) );
BUF_X1 \mylsu/_2459_ ( .A(\mylsu/araddr_tmp [9] ), .Z(\mylsu/_0077_ ) );
BUF_X1 \mylsu/_2460_ ( .A(\EX_LS_dest_csreg_mem [9] ), .Z(\mylsu/_0341_ ) );
BUF_X1 \mylsu/_2461_ ( .A(\mylsu/_0045_ ), .Z(\araddr_LSU [9] ) );
BUF_X1 \mylsu/_2462_ ( .A(\mylsu/araddr_tmp [10] ), .Z(\mylsu/_0047_ ) );
BUF_X1 \mylsu/_2463_ ( .A(\EX_LS_dest_csreg_mem [10] ), .Z(\mylsu/_0311_ ) );
BUF_X1 \mylsu/_2464_ ( .A(\mylsu/_0015_ ), .Z(\araddr_LSU [10] ) );
BUF_X1 \mylsu/_2465_ ( .A(\mylsu/araddr_tmp [11] ), .Z(\mylsu/_0048_ ) );
BUF_X1 \mylsu/_2466_ ( .A(\EX_LS_dest_csreg_mem [11] ), .Z(\mylsu/_0312_ ) );
BUF_X1 \mylsu/_2467_ ( .A(\mylsu/_0016_ ), .Z(\araddr_LSU [11] ) );
BUF_X1 \mylsu/_2468_ ( .A(\mylsu/araddr_tmp [12] ), .Z(\mylsu/_0049_ ) );
BUF_X1 \mylsu/_2469_ ( .A(\EX_LS_dest_csreg_mem [12] ), .Z(\mylsu/_0313_ ) );
BUF_X1 \mylsu/_2470_ ( .A(\mylsu/_0017_ ), .Z(\araddr_LSU [12] ) );
BUF_X1 \mylsu/_2471_ ( .A(\mylsu/araddr_tmp [13] ), .Z(\mylsu/_0050_ ) );
BUF_X1 \mylsu/_2472_ ( .A(\EX_LS_dest_csreg_mem [13] ), .Z(\mylsu/_0314_ ) );
BUF_X1 \mylsu/_2473_ ( .A(\mylsu/_0018_ ), .Z(\araddr_LSU [13] ) );
BUF_X1 \mylsu/_2474_ ( .A(\mylsu/araddr_tmp [14] ), .Z(\mylsu/_0051_ ) );
BUF_X1 \mylsu/_2475_ ( .A(\EX_LS_dest_csreg_mem [14] ), .Z(\mylsu/_0315_ ) );
BUF_X1 \mylsu/_2476_ ( .A(\mylsu/_0019_ ), .Z(\araddr_LSU [14] ) );
BUF_X1 \mylsu/_2477_ ( .A(\mylsu/araddr_tmp [15] ), .Z(\mylsu/_0052_ ) );
BUF_X1 \mylsu/_2478_ ( .A(\EX_LS_dest_csreg_mem [15] ), .Z(\mylsu/_0316_ ) );
BUF_X1 \mylsu/_2479_ ( .A(\mylsu/_0020_ ), .Z(\araddr_LSU [15] ) );
BUF_X1 \mylsu/_2480_ ( .A(\mylsu/araddr_tmp [16] ), .Z(\mylsu/_0053_ ) );
BUF_X1 \mylsu/_2481_ ( .A(\EX_LS_dest_csreg_mem [16] ), .Z(\mylsu/_0317_ ) );
BUF_X1 \mylsu/_2482_ ( .A(\mylsu/_0021_ ), .Z(\araddr_LSU [16] ) );
BUF_X1 \mylsu/_2483_ ( .A(\mylsu/araddr_tmp [17] ), .Z(\mylsu/_0054_ ) );
BUF_X1 \mylsu/_2484_ ( .A(\EX_LS_dest_csreg_mem [17] ), .Z(\mylsu/_0318_ ) );
BUF_X1 \mylsu/_2485_ ( .A(\mylsu/_0022_ ), .Z(\araddr_LSU [17] ) );
BUF_X1 \mylsu/_2486_ ( .A(\mylsu/araddr_tmp [18] ), .Z(\mylsu/_0055_ ) );
BUF_X1 \mylsu/_2487_ ( .A(\EX_LS_dest_csreg_mem [18] ), .Z(\mylsu/_0319_ ) );
BUF_X1 \mylsu/_2488_ ( .A(\mylsu/_0023_ ), .Z(\araddr_LSU [18] ) );
BUF_X1 \mylsu/_2489_ ( .A(\mylsu/araddr_tmp [19] ), .Z(\mylsu/_0056_ ) );
BUF_X1 \mylsu/_2490_ ( .A(\EX_LS_dest_csreg_mem [19] ), .Z(\mylsu/_0320_ ) );
BUF_X1 \mylsu/_2491_ ( .A(\mylsu/_0024_ ), .Z(\araddr_LSU [19] ) );
BUF_X1 \mylsu/_2492_ ( .A(\mylsu/araddr_tmp [20] ), .Z(\mylsu/_0058_ ) );
BUF_X1 \mylsu/_2493_ ( .A(\EX_LS_dest_csreg_mem [20] ), .Z(\mylsu/_0322_ ) );
BUF_X1 \mylsu/_2494_ ( .A(\mylsu/_0026_ ), .Z(\araddr_LSU [20] ) );
BUF_X1 \mylsu/_2495_ ( .A(\mylsu/araddr_tmp [21] ), .Z(\mylsu/_0059_ ) );
BUF_X1 \mylsu/_2496_ ( .A(\EX_LS_dest_csreg_mem [21] ), .Z(\mylsu/_0323_ ) );
BUF_X1 \mylsu/_2497_ ( .A(\mylsu/_0027_ ), .Z(\araddr_LSU [21] ) );
BUF_X1 \mylsu/_2498_ ( .A(\mylsu/araddr_tmp [22] ), .Z(\mylsu/_0060_ ) );
BUF_X1 \mylsu/_2499_ ( .A(\EX_LS_dest_csreg_mem [22] ), .Z(\mylsu/_0324_ ) );
BUF_X1 \mylsu/_2500_ ( .A(\mylsu/_0028_ ), .Z(\araddr_LSU [22] ) );
BUF_X1 \mylsu/_2501_ ( .A(\mylsu/araddr_tmp [23] ), .Z(\mylsu/_0061_ ) );
BUF_X1 \mylsu/_2502_ ( .A(\EX_LS_dest_csreg_mem [23] ), .Z(\mylsu/_0325_ ) );
BUF_X1 \mylsu/_2503_ ( .A(\mylsu/_0029_ ), .Z(\araddr_LSU [23] ) );
BUF_X1 \mylsu/_2504_ ( .A(\mylsu/araddr_tmp [24] ), .Z(\mylsu/_0062_ ) );
BUF_X1 \mylsu/_2505_ ( .A(\EX_LS_dest_csreg_mem [24] ), .Z(\mylsu/_0326_ ) );
BUF_X1 \mylsu/_2506_ ( .A(\mylsu/_0030_ ), .Z(\araddr_LSU [24] ) );
BUF_X1 \mylsu/_2507_ ( .A(\mylsu/araddr_tmp [25] ), .Z(\mylsu/_0063_ ) );
BUF_X1 \mylsu/_2508_ ( .A(\EX_LS_dest_csreg_mem [25] ), .Z(\mylsu/_0327_ ) );
BUF_X1 \mylsu/_2509_ ( .A(\mylsu/_0031_ ), .Z(\araddr_LSU [25] ) );
BUF_X1 \mylsu/_2510_ ( .A(\mylsu/araddr_tmp [26] ), .Z(\mylsu/_0064_ ) );
BUF_X1 \mylsu/_2511_ ( .A(\EX_LS_dest_csreg_mem [26] ), .Z(\mylsu/_0328_ ) );
BUF_X1 \mylsu/_2512_ ( .A(\mylsu/_0032_ ), .Z(\araddr_LSU [26] ) );
BUF_X1 \mylsu/_2513_ ( .A(\mylsu/araddr_tmp [27] ), .Z(\mylsu/_0065_ ) );
BUF_X1 \mylsu/_2514_ ( .A(\EX_LS_dest_csreg_mem [27] ), .Z(\mylsu/_0329_ ) );
BUF_X1 \mylsu/_2515_ ( .A(\mylsu/_0033_ ), .Z(\araddr_LSU [27] ) );
BUF_X1 \mylsu/_2516_ ( .A(\mylsu/araddr_tmp [28] ), .Z(\mylsu/_0066_ ) );
BUF_X1 \mylsu/_2517_ ( .A(\EX_LS_dest_csreg_mem [28] ), .Z(\mylsu/_0330_ ) );
BUF_X1 \mylsu/_2518_ ( .A(\mylsu/_0034_ ), .Z(\araddr_LSU [28] ) );
BUF_X1 \mylsu/_2519_ ( .A(\mylsu/araddr_tmp [29] ), .Z(\mylsu/_0067_ ) );
BUF_X1 \mylsu/_2520_ ( .A(\EX_LS_dest_csreg_mem [29] ), .Z(\mylsu/_0331_ ) );
BUF_X1 \mylsu/_2521_ ( .A(\mylsu/_0035_ ), .Z(\araddr_LSU [29] ) );
BUF_X1 \mylsu/_2522_ ( .A(\mylsu/araddr_tmp [30] ), .Z(\mylsu/_0069_ ) );
BUF_X1 \mylsu/_2523_ ( .A(\EX_LS_dest_csreg_mem [30] ), .Z(\mylsu/_0333_ ) );
BUF_X1 \mylsu/_2524_ ( .A(\mylsu/_0037_ ), .Z(\araddr_LSU [30] ) );
BUF_X1 \mylsu/_2525_ ( .A(\mylsu/araddr_tmp [31] ), .Z(\mylsu/_0070_ ) );
BUF_X1 \mylsu/_2526_ ( .A(\EX_LS_dest_csreg_mem [31] ), .Z(\mylsu/_0334_ ) );
BUF_X1 \mylsu/_2527_ ( .A(\mylsu/_0038_ ), .Z(\araddr_LSU [31] ) );
BUF_X1 \mylsu/_2528_ ( .A(\EX_LS_typ [1] ), .Z(\mylsu/_0919_ ) );
BUF_X1 \mylsu/_2529_ ( .A(\EX_LS_typ [0] ), .Z(\mylsu/_0918_ ) );
BUF_X1 \mylsu/_2530_ ( .A(\EX_LS_typ [3] ), .Z(\mylsu/_0921_ ) );
BUF_X1 \mylsu/_2531_ ( .A(\EX_LS_typ [2] ), .Z(\mylsu/_0920_ ) );
BUF_X1 \mylsu/_2532_ ( .A(\EX_LS_typ [4] ), .Z(\mylsu/_0922_ ) );
BUF_X1 \mylsu/_2533_ ( .A(\mylsu/_0299_ ), .Z(\awsize_LSU [0] ) );
BUF_X1 \mylsu/_2534_ ( .A(\mylsu/_0300_ ), .Z(\awsize_LSU [1] ) );
BUF_X1 \mylsu/_2535_ ( .A(\mylsu/awaddr_tmp [0] ), .Z(\mylsu/_0266_ ) );
BUF_X1 \mylsu/_2536_ ( .A(\mylsu/_0234_ ), .Z(\awaddr_LSU [0] ) );
BUF_X1 \mylsu/_2537_ ( .A(\mylsu/awaddr_tmp [1] ), .Z(\mylsu/_0277_ ) );
BUF_X1 \mylsu/_2538_ ( .A(\mylsu/_0245_ ), .Z(\awaddr_LSU [1] ) );
BUF_X1 \mylsu/_2539_ ( .A(\mylsu/awaddr_tmp [2] ), .Z(\mylsu/_0288_ ) );
BUF_X1 \mylsu/_2540_ ( .A(\mylsu/_0256_ ), .Z(\awaddr_LSU [2] ) );
BUF_X1 \mylsu/_2541_ ( .A(\mylsu/awaddr_tmp [3] ), .Z(\mylsu/_0291_ ) );
BUF_X1 \mylsu/_2542_ ( .A(\mylsu/_0259_ ), .Z(\awaddr_LSU [3] ) );
BUF_X1 \mylsu/_2543_ ( .A(\mylsu/awaddr_tmp [4] ), .Z(\mylsu/_0292_ ) );
BUF_X1 \mylsu/_2544_ ( .A(\mylsu/_0260_ ), .Z(\awaddr_LSU [4] ) );
BUF_X1 \mylsu/_2545_ ( .A(\mylsu/awaddr_tmp [5] ), .Z(\mylsu/_0293_ ) );
BUF_X1 \mylsu/_2546_ ( .A(\mylsu/_0261_ ), .Z(\awaddr_LSU [5] ) );
BUF_X1 \mylsu/_2547_ ( .A(\mylsu/awaddr_tmp [6] ), .Z(\mylsu/_0294_ ) );
BUF_X1 \mylsu/_2548_ ( .A(\mylsu/_0262_ ), .Z(\awaddr_LSU [6] ) );
BUF_X1 \mylsu/_2549_ ( .A(\mylsu/awaddr_tmp [7] ), .Z(\mylsu/_0295_ ) );
BUF_X1 \mylsu/_2550_ ( .A(\mylsu/_0263_ ), .Z(\awaddr_LSU [7] ) );
BUF_X1 \mylsu/_2551_ ( .A(\mylsu/awaddr_tmp [8] ), .Z(\mylsu/_0296_ ) );
BUF_X1 \mylsu/_2552_ ( .A(\mylsu/_0264_ ), .Z(\awaddr_LSU [8] ) );
BUF_X1 \mylsu/_2553_ ( .A(\mylsu/awaddr_tmp [9] ), .Z(\mylsu/_0297_ ) );
BUF_X1 \mylsu/_2554_ ( .A(\mylsu/_0265_ ), .Z(\awaddr_LSU [9] ) );
BUF_X1 \mylsu/_2555_ ( .A(\mylsu/awaddr_tmp [10] ), .Z(\mylsu/_0267_ ) );
BUF_X1 \mylsu/_2556_ ( .A(\mylsu/_0235_ ), .Z(\awaddr_LSU [10] ) );
BUF_X1 \mylsu/_2557_ ( .A(\mylsu/awaddr_tmp [11] ), .Z(\mylsu/_0268_ ) );
BUF_X1 \mylsu/_2558_ ( .A(\mylsu/_0236_ ), .Z(\awaddr_LSU [11] ) );
BUF_X1 \mylsu/_2559_ ( .A(\mylsu/awaddr_tmp [12] ), .Z(\mylsu/_0269_ ) );
BUF_X1 \mylsu/_2560_ ( .A(\mylsu/_0237_ ), .Z(\awaddr_LSU [12] ) );
BUF_X1 \mylsu/_2561_ ( .A(\mylsu/awaddr_tmp [13] ), .Z(\mylsu/_0270_ ) );
BUF_X1 \mylsu/_2562_ ( .A(\mylsu/_0238_ ), .Z(\awaddr_LSU [13] ) );
BUF_X1 \mylsu/_2563_ ( .A(\mylsu/awaddr_tmp [14] ), .Z(\mylsu/_0271_ ) );
BUF_X1 \mylsu/_2564_ ( .A(\mylsu/_0239_ ), .Z(\awaddr_LSU [14] ) );
BUF_X1 \mylsu/_2565_ ( .A(\mylsu/awaddr_tmp [15] ), .Z(\mylsu/_0272_ ) );
BUF_X1 \mylsu/_2566_ ( .A(\mylsu/_0240_ ), .Z(\awaddr_LSU [15] ) );
BUF_X1 \mylsu/_2567_ ( .A(\mylsu/awaddr_tmp [16] ), .Z(\mylsu/_0273_ ) );
BUF_X1 \mylsu/_2568_ ( .A(\mylsu/_0241_ ), .Z(\awaddr_LSU [16] ) );
BUF_X1 \mylsu/_2569_ ( .A(\mylsu/awaddr_tmp [17] ), .Z(\mylsu/_0274_ ) );
BUF_X1 \mylsu/_2570_ ( .A(\mylsu/_0242_ ), .Z(\awaddr_LSU [17] ) );
BUF_X1 \mylsu/_2571_ ( .A(\mylsu/awaddr_tmp [18] ), .Z(\mylsu/_0275_ ) );
BUF_X1 \mylsu/_2572_ ( .A(\mylsu/_0243_ ), .Z(\awaddr_LSU [18] ) );
BUF_X1 \mylsu/_2573_ ( .A(\mylsu/awaddr_tmp [19] ), .Z(\mylsu/_0276_ ) );
BUF_X1 \mylsu/_2574_ ( .A(\mylsu/_0244_ ), .Z(\awaddr_LSU [19] ) );
BUF_X1 \mylsu/_2575_ ( .A(\mylsu/awaddr_tmp [20] ), .Z(\mylsu/_0278_ ) );
BUF_X1 \mylsu/_2576_ ( .A(\mylsu/_0246_ ), .Z(\awaddr_LSU [20] ) );
BUF_X1 \mylsu/_2577_ ( .A(\mylsu/awaddr_tmp [21] ), .Z(\mylsu/_0279_ ) );
BUF_X1 \mylsu/_2578_ ( .A(\mylsu/_0247_ ), .Z(\awaddr_LSU [21] ) );
BUF_X1 \mylsu/_2579_ ( .A(\mylsu/awaddr_tmp [22] ), .Z(\mylsu/_0280_ ) );
BUF_X1 \mylsu/_2580_ ( .A(\mylsu/_0248_ ), .Z(\awaddr_LSU [22] ) );
BUF_X1 \mylsu/_2581_ ( .A(\mylsu/awaddr_tmp [23] ), .Z(\mylsu/_0281_ ) );
BUF_X1 \mylsu/_2582_ ( .A(\mylsu/_0249_ ), .Z(\awaddr_LSU [23] ) );
BUF_X1 \mylsu/_2583_ ( .A(\mylsu/awaddr_tmp [24] ), .Z(\mylsu/_0282_ ) );
BUF_X1 \mylsu/_2584_ ( .A(\mylsu/_0250_ ), .Z(\awaddr_LSU [24] ) );
BUF_X1 \mylsu/_2585_ ( .A(\mylsu/awaddr_tmp [25] ), .Z(\mylsu/_0283_ ) );
BUF_X1 \mylsu/_2586_ ( .A(\mylsu/_0251_ ), .Z(\awaddr_LSU [25] ) );
BUF_X1 \mylsu/_2587_ ( .A(\mylsu/awaddr_tmp [26] ), .Z(\mylsu/_0284_ ) );
BUF_X1 \mylsu/_2588_ ( .A(\mylsu/_0252_ ), .Z(\awaddr_LSU [26] ) );
BUF_X1 \mylsu/_2589_ ( .A(\mylsu/awaddr_tmp [27] ), .Z(\mylsu/_0285_ ) );
BUF_X1 \mylsu/_2590_ ( .A(\mylsu/_0253_ ), .Z(\awaddr_LSU [27] ) );
BUF_X1 \mylsu/_2591_ ( .A(\mylsu/awaddr_tmp [28] ), .Z(\mylsu/_0286_ ) );
BUF_X1 \mylsu/_2592_ ( .A(\mylsu/_0254_ ), .Z(\awaddr_LSU [28] ) );
BUF_X1 \mylsu/_2593_ ( .A(\mylsu/awaddr_tmp [29] ), .Z(\mylsu/_0287_ ) );
BUF_X1 \mylsu/_2594_ ( .A(\mylsu/_0255_ ), .Z(\awaddr_LSU [29] ) );
BUF_X1 \mylsu/_2595_ ( .A(\mylsu/awaddr_tmp [30] ), .Z(\mylsu/_0289_ ) );
BUF_X1 \mylsu/_2596_ ( .A(\mylsu/_0257_ ), .Z(\awaddr_LSU [30] ) );
BUF_X1 \mylsu/_2597_ ( .A(\mylsu/awaddr_tmp [31] ), .Z(\mylsu/_0290_ ) );
BUF_X1 \mylsu/_2598_ ( .A(\mylsu/_0258_ ), .Z(\awaddr_LSU [31] ) );
BUF_X1 \mylsu/_2599_ ( .A(\mylsu/_0947_ ), .Z(\wdata_LSU [0] ) );
BUF_X1 \mylsu/_2600_ ( .A(\mylsu/_0958_ ), .Z(\wdata_LSU [1] ) );
BUF_X1 \mylsu/_2601_ ( .A(\mylsu/_0969_ ), .Z(\wdata_LSU [2] ) );
BUF_X1 \mylsu/_2602_ ( .A(\mylsu/_0972_ ), .Z(\wdata_LSU [3] ) );
BUF_X1 \mylsu/_2603_ ( .A(\mylsu/_0973_ ), .Z(\wdata_LSU [4] ) );
BUF_X1 \mylsu/_2604_ ( .A(\mylsu/_0974_ ), .Z(\wdata_LSU [5] ) );
BUF_X1 \mylsu/_2605_ ( .A(\mylsu/_0975_ ), .Z(\wdata_LSU [6] ) );
BUF_X1 \mylsu/_2606_ ( .A(\mylsu/_0976_ ), .Z(\wdata_LSU [7] ) );
BUF_X1 \mylsu/_2607_ ( .A(\mylsu/_0977_ ), .Z(\wdata_LSU [8] ) );
BUF_X1 \mylsu/_2608_ ( .A(\mylsu/_0978_ ), .Z(\wdata_LSU [9] ) );
BUF_X1 \mylsu/_2609_ ( .A(\mylsu/_0948_ ), .Z(\wdata_LSU [10] ) );
BUF_X1 \mylsu/_2610_ ( .A(\mylsu/_0949_ ), .Z(\wdata_LSU [11] ) );
BUF_X1 \mylsu/_2611_ ( .A(\mylsu/_0950_ ), .Z(\wdata_LSU [12] ) );
BUF_X1 \mylsu/_2612_ ( .A(\mylsu/_0951_ ), .Z(\wdata_LSU [13] ) );
BUF_X1 \mylsu/_2613_ ( .A(\mylsu/_0952_ ), .Z(\wdata_LSU [14] ) );
BUF_X1 \mylsu/_2614_ ( .A(\mylsu/_0953_ ), .Z(\wdata_LSU [15] ) );
BUF_X1 \mylsu/_2615_ ( .A(\mylsu/_0954_ ), .Z(\wdata_LSU [16] ) );
BUF_X1 \mylsu/_2616_ ( .A(\mylsu/_0955_ ), .Z(\wdata_LSU [17] ) );
BUF_X1 \mylsu/_2617_ ( .A(\mylsu/_0956_ ), .Z(\wdata_LSU [18] ) );
BUF_X1 \mylsu/_2618_ ( .A(\mylsu/_0957_ ), .Z(\wdata_LSU [19] ) );
BUF_X1 \mylsu/_2619_ ( .A(\mylsu/_0959_ ), .Z(\wdata_LSU [20] ) );
BUF_X1 \mylsu/_2620_ ( .A(\mylsu/_0960_ ), .Z(\wdata_LSU [21] ) );
BUF_X1 \mylsu/_2621_ ( .A(\mylsu/_0961_ ), .Z(\wdata_LSU [22] ) );
BUF_X1 \mylsu/_2622_ ( .A(\mylsu/_0962_ ), .Z(\wdata_LSU [23] ) );
BUF_X1 \mylsu/_2623_ ( .A(\mylsu/_0963_ ), .Z(\wdata_LSU [24] ) );
BUF_X1 \mylsu/_2624_ ( .A(\mylsu/_0964_ ), .Z(\wdata_LSU [25] ) );
BUF_X1 \mylsu/_2625_ ( .A(\mylsu/_0965_ ), .Z(\wdata_LSU [26] ) );
BUF_X1 \mylsu/_2626_ ( .A(\mylsu/_0966_ ), .Z(\wdata_LSU [27] ) );
BUF_X1 \mylsu/_2627_ ( .A(\mylsu/_0967_ ), .Z(\wdata_LSU [28] ) );
BUF_X1 \mylsu/_2628_ ( .A(\mylsu/_0968_ ), .Z(\wdata_LSU [29] ) );
BUF_X1 \mylsu/_2629_ ( .A(\mylsu/_0970_ ), .Z(\wdata_LSU [30] ) );
BUF_X1 \mylsu/_2630_ ( .A(\mylsu/_0971_ ), .Z(\wdata_LSU [31] ) );
BUF_X1 \mylsu/_2631_ ( .A(\mylsu/_1048_ ), .Z(\wstrb_LSU [0] ) );
BUF_X1 \mylsu/_2632_ ( .A(\mylsu/_1049_ ), .Z(\wstrb_LSU [1] ) );
BUF_X1 \mylsu/_2633_ ( .A(\mylsu/_1050_ ), .Z(\wstrb_LSU [2] ) );
BUF_X1 \mylsu/_2634_ ( .A(\mylsu/_1051_ ), .Z(\wstrb_LSU [3] ) );
BUF_X1 \mylsu/_2635_ ( .A(LS_WB_pc ), .Z(\mylsu/_0804_ ) );
BUF_X1 \mylsu/_2636_ ( .A(\LS_WB_waddr_reg [0] ), .Z(\mylsu/_0942_ ) );
BUF_X1 \mylsu/_2637_ ( .A(\EX_LS_dest_reg [0] ), .Z(\mylsu/_0342_ ) );
BUF_X1 \mylsu/_2638_ ( .A(\mylsu/_0081_ ), .Z(\mylsu/_1213_ ) );
BUF_X1 \mylsu/_2639_ ( .A(\LS_WB_waddr_reg [1] ), .Z(\mylsu/_0943_ ) );
BUF_X1 \mylsu/_2640_ ( .A(\EX_LS_dest_reg [1] ), .Z(\mylsu/_0343_ ) );
BUF_X1 \mylsu/_2641_ ( .A(\mylsu/_0082_ ), .Z(\mylsu/_1214_ ) );
BUF_X1 \mylsu/_2642_ ( .A(\LS_WB_waddr_reg [2] ), .Z(\mylsu/_0944_ ) );
BUF_X1 \mylsu/_2643_ ( .A(\EX_LS_dest_reg [2] ), .Z(\mylsu/_0344_ ) );
BUF_X1 \mylsu/_2644_ ( .A(\mylsu/_0083_ ), .Z(\mylsu/_1215_ ) );
BUF_X1 \mylsu/_2645_ ( .A(\LS_WB_waddr_reg [3] ), .Z(\mylsu/_0945_ ) );
BUF_X1 \mylsu/_2646_ ( .A(\EX_LS_dest_reg [3] ), .Z(\mylsu/_0345_ ) );
BUF_X1 \mylsu/_2647_ ( .A(\mylsu/_0084_ ), .Z(\mylsu/_1216_ ) );
BUF_X1 \mylsu/_2648_ ( .A(\LS_WB_waddr_reg [4] ), .Z(\mylsu/_0946_ ) );
BUF_X1 \mylsu/_2649_ ( .A(\EX_LS_dest_reg [4] ), .Z(\mylsu/_0346_ ) );
BUF_X1 \mylsu/_2650_ ( .A(\mylsu/_0085_ ), .Z(\mylsu/_1217_ ) );
BUF_X1 \mylsu/_2651_ ( .A(\LS_WB_waddr_csreg [0] ), .Z(\mylsu/_0930_ ) );
BUF_X1 \mylsu/_2652_ ( .A(\mylsu/_0086_ ), .Z(\mylsu/_1218_ ) );
BUF_X1 \mylsu/_2653_ ( .A(\LS_WB_waddr_csreg [1] ), .Z(\mylsu/_0933_ ) );
BUF_X1 \mylsu/_2654_ ( .A(\mylsu/_0087_ ), .Z(\mylsu/_1219_ ) );
BUF_X1 \mylsu/_2655_ ( .A(\LS_WB_waddr_csreg [2] ), .Z(\mylsu/_0934_ ) );
BUF_X1 \mylsu/_2656_ ( .A(\mylsu/_0088_ ), .Z(\mylsu/_1220_ ) );
BUF_X1 \mylsu/_2657_ ( .A(\LS_WB_waddr_csreg [3] ), .Z(\mylsu/_0935_ ) );
BUF_X1 \mylsu/_2658_ ( .A(\mylsu/_0089_ ), .Z(\mylsu/_1221_ ) );
BUF_X1 \mylsu/_2659_ ( .A(\LS_WB_waddr_csreg [4] ), .Z(\mylsu/_0936_ ) );
BUF_X1 \mylsu/_2660_ ( .A(\mylsu/_0090_ ), .Z(\mylsu/_1222_ ) );
BUF_X1 \mylsu/_2661_ ( .A(\LS_WB_waddr_csreg [5] ), .Z(\mylsu/_0937_ ) );
BUF_X1 \mylsu/_2662_ ( .A(\mylsu/_0091_ ), .Z(\mylsu/_1223_ ) );
BUF_X1 \mylsu/_2663_ ( .A(\LS_WB_waddr_csreg [6] ), .Z(\mylsu/_0938_ ) );
BUF_X1 \mylsu/_2664_ ( .A(\mylsu/_0092_ ), .Z(\mylsu/_1224_ ) );
BUF_X1 \mylsu/_2665_ ( .A(\LS_WB_waddr_csreg [7] ), .Z(\mylsu/_0939_ ) );
BUF_X1 \mylsu/_2666_ ( .A(\mylsu/_0093_ ), .Z(\mylsu/_1225_ ) );
BUF_X1 \mylsu/_2667_ ( .A(\LS_WB_waddr_csreg [8] ), .Z(\mylsu/_0940_ ) );
BUF_X1 \mylsu/_2668_ ( .A(\mylsu/_0094_ ), .Z(\mylsu/_1226_ ) );
BUF_X1 \mylsu/_2669_ ( .A(\LS_WB_waddr_csreg [9] ), .Z(\mylsu/_0941_ ) );
BUF_X1 \mylsu/_2670_ ( .A(\mylsu/_0095_ ), .Z(\mylsu/_1227_ ) );
BUF_X1 \mylsu/_2671_ ( .A(\LS_WB_waddr_csreg [10] ), .Z(\mylsu/_0931_ ) );
BUF_X1 \mylsu/_2672_ ( .A(\mylsu/_0096_ ), .Z(\mylsu/_1228_ ) );
BUF_X1 \mylsu/_2673_ ( .A(\LS_WB_waddr_csreg [11] ), .Z(\mylsu/_0932_ ) );
BUF_X1 \mylsu/_2674_ ( .A(\mylsu/_0097_ ), .Z(\mylsu/_1229_ ) );
BUF_X1 \mylsu/_2675_ ( .A(\LS_WB_wdata_reg [0] ), .Z(\mylsu/_1011_ ) );
BUF_X1 \mylsu/_2676_ ( .A(\mylsu/_0098_ ), .Z(\mylsu/_1230_ ) );
BUF_X1 \mylsu/_2677_ ( .A(\LS_WB_wdata_reg [1] ), .Z(\mylsu/_1022_ ) );
BUF_X1 \mylsu/_2678_ ( .A(\mylsu/_0099_ ), .Z(\mylsu/_1231_ ) );
BUF_X1 \mylsu/_2679_ ( .A(\LS_WB_wdata_reg [2] ), .Z(\mylsu/_1033_ ) );
BUF_X1 \mylsu/_2680_ ( .A(\mylsu/_0100_ ), .Z(\mylsu/_1232_ ) );
BUF_X1 \mylsu/_2681_ ( .A(\LS_WB_wdata_reg [3] ), .Z(\mylsu/_1036_ ) );
BUF_X1 \mylsu/_2682_ ( .A(\mylsu/_0101_ ), .Z(\mylsu/_1233_ ) );
BUF_X1 \mylsu/_2683_ ( .A(\LS_WB_wdata_reg [4] ), .Z(\mylsu/_1037_ ) );
BUF_X1 \mylsu/_2684_ ( .A(\mylsu/_0102_ ), .Z(\mylsu/_1234_ ) );
BUF_X1 \mylsu/_2685_ ( .A(\LS_WB_wdata_reg [5] ), .Z(\mylsu/_1038_ ) );
BUF_X1 \mylsu/_2686_ ( .A(\mylsu/_0103_ ), .Z(\mylsu/_1235_ ) );
BUF_X1 \mylsu/_2687_ ( .A(\LS_WB_wdata_reg [6] ), .Z(\mylsu/_1039_ ) );
BUF_X1 \mylsu/_2688_ ( .A(\mylsu/_0104_ ), .Z(\mylsu/_1236_ ) );
BUF_X1 \mylsu/_2689_ ( .A(\LS_WB_wdata_reg [7] ), .Z(\mylsu/_1040_ ) );
BUF_X1 \mylsu/_2690_ ( .A(\mylsu/_0105_ ), .Z(\mylsu/_1237_ ) );
BUF_X1 \mylsu/_2691_ ( .A(\LS_WB_wdata_reg [8] ), .Z(\mylsu/_1041_ ) );
BUF_X1 \mylsu/_2692_ ( .A(\mylsu/_0106_ ), .Z(\mylsu/_1238_ ) );
BUF_X1 \mylsu/_2693_ ( .A(\LS_WB_wdata_reg [9] ), .Z(\mylsu/_1042_ ) );
BUF_X1 \mylsu/_2694_ ( .A(\mylsu/_0107_ ), .Z(\mylsu/_1239_ ) );
BUF_X1 \mylsu/_2695_ ( .A(\LS_WB_wdata_reg [10] ), .Z(\mylsu/_1012_ ) );
BUF_X1 \mylsu/_2696_ ( .A(\mylsu/_0108_ ), .Z(\mylsu/_1240_ ) );
BUF_X1 \mylsu/_2697_ ( .A(\LS_WB_wdata_reg [11] ), .Z(\mylsu/_1013_ ) );
BUF_X1 \mylsu/_2698_ ( .A(\mylsu/_0109_ ), .Z(\mylsu/_1241_ ) );
BUF_X1 \mylsu/_2699_ ( .A(\LS_WB_wdata_reg [12] ), .Z(\mylsu/_1014_ ) );
BUF_X1 \mylsu/_2700_ ( .A(\mylsu/_0110_ ), .Z(\mylsu/_1242_ ) );
BUF_X1 \mylsu/_2701_ ( .A(\LS_WB_wdata_reg [13] ), .Z(\mylsu/_1015_ ) );
BUF_X1 \mylsu/_2702_ ( .A(\mylsu/_0111_ ), .Z(\mylsu/_1243_ ) );
BUF_X1 \mylsu/_2703_ ( .A(\LS_WB_wdata_reg [14] ), .Z(\mylsu/_1016_ ) );
BUF_X1 \mylsu/_2704_ ( .A(\mylsu/_0112_ ), .Z(\mylsu/_1244_ ) );
BUF_X1 \mylsu/_2705_ ( .A(\LS_WB_wdata_reg [15] ), .Z(\mylsu/_1017_ ) );
BUF_X1 \mylsu/_2706_ ( .A(\mylsu/_0113_ ), .Z(\mylsu/_1245_ ) );
BUF_X1 \mylsu/_2707_ ( .A(\LS_WB_wdata_reg [16] ), .Z(\mylsu/_1018_ ) );
BUF_X1 \mylsu/_2708_ ( .A(\mylsu/_0114_ ), .Z(\mylsu/_1246_ ) );
BUF_X1 \mylsu/_2709_ ( .A(\LS_WB_wdata_reg [17] ), .Z(\mylsu/_1019_ ) );
BUF_X1 \mylsu/_2710_ ( .A(\mylsu/_0115_ ), .Z(\mylsu/_1247_ ) );
BUF_X1 \mylsu/_2711_ ( .A(\LS_WB_wdata_reg [18] ), .Z(\mylsu/_1020_ ) );
BUF_X1 \mylsu/_2712_ ( .A(\mylsu/_0116_ ), .Z(\mylsu/_1248_ ) );
BUF_X1 \mylsu/_2713_ ( .A(\LS_WB_wdata_reg [19] ), .Z(\mylsu/_1021_ ) );
BUF_X1 \mylsu/_2714_ ( .A(\mylsu/_0117_ ), .Z(\mylsu/_1249_ ) );
BUF_X1 \mylsu/_2715_ ( .A(\LS_WB_wdata_reg [20] ), .Z(\mylsu/_1023_ ) );
BUF_X1 \mylsu/_2716_ ( .A(\mylsu/_0118_ ), .Z(\mylsu/_1250_ ) );
BUF_X1 \mylsu/_2717_ ( .A(\LS_WB_wdata_reg [21] ), .Z(\mylsu/_1024_ ) );
BUF_X1 \mylsu/_2718_ ( .A(\mylsu/_0119_ ), .Z(\mylsu/_1251_ ) );
BUF_X1 \mylsu/_2719_ ( .A(\LS_WB_wdata_reg [22] ), .Z(\mylsu/_1025_ ) );
BUF_X1 \mylsu/_2720_ ( .A(\mylsu/_0120_ ), .Z(\mylsu/_1252_ ) );
BUF_X1 \mylsu/_2721_ ( .A(\LS_WB_wdata_reg [23] ), .Z(\mylsu/_1026_ ) );
BUF_X1 \mylsu/_2722_ ( .A(\mylsu/_0121_ ), .Z(\mylsu/_1253_ ) );
BUF_X1 \mylsu/_2723_ ( .A(\LS_WB_wdata_reg [24] ), .Z(\mylsu/_1027_ ) );
BUF_X1 \mylsu/_2724_ ( .A(\mylsu/_0122_ ), .Z(\mylsu/_1254_ ) );
BUF_X1 \mylsu/_2725_ ( .A(\LS_WB_wdata_reg [25] ), .Z(\mylsu/_1028_ ) );
BUF_X1 \mylsu/_2726_ ( .A(\mylsu/_0123_ ), .Z(\mylsu/_1255_ ) );
BUF_X1 \mylsu/_2727_ ( .A(\LS_WB_wdata_reg [26] ), .Z(\mylsu/_1029_ ) );
BUF_X1 \mylsu/_2728_ ( .A(\mylsu/_0124_ ), .Z(\mylsu/_1256_ ) );
BUF_X1 \mylsu/_2729_ ( .A(\LS_WB_wdata_reg [27] ), .Z(\mylsu/_1030_ ) );
BUF_X1 \mylsu/_2730_ ( .A(\mylsu/_0125_ ), .Z(\mylsu/_1257_ ) );
BUF_X1 \mylsu/_2731_ ( .A(\LS_WB_wdata_reg [28] ), .Z(\mylsu/_1031_ ) );
BUF_X1 \mylsu/_2732_ ( .A(\mylsu/_0126_ ), .Z(\mylsu/_1258_ ) );
BUF_X1 \mylsu/_2733_ ( .A(\LS_WB_wdata_reg [29] ), .Z(\mylsu/_1032_ ) );
BUF_X1 \mylsu/_2734_ ( .A(\mylsu/_0127_ ), .Z(\mylsu/_1259_ ) );
BUF_X1 \mylsu/_2735_ ( .A(\LS_WB_wdata_reg [30] ), .Z(\mylsu/_1034_ ) );
BUF_X1 \mylsu/_2736_ ( .A(\mylsu/_0128_ ), .Z(\mylsu/_1260_ ) );
BUF_X1 \mylsu/_2737_ ( .A(\LS_WB_wdata_reg [31] ), .Z(\mylsu/_1035_ ) );
BUF_X1 \mylsu/_2738_ ( .A(\mylsu/_0129_ ), .Z(\mylsu/_1261_ ) );
BUF_X1 \mylsu/_2739_ ( .A(LS_WB_wen_reg ), .Z(\mylsu/_1046_ ) );
BUF_X1 \mylsu/_2740_ ( .A(previous_load_done ), .Z(\mylsu/_0805_ ) );
BUF_X1 \mylsu/_2741_ ( .A(\LS_WB_wdata_csreg [0] ), .Z(\mylsu/_0979_ ) );
BUF_X1 \mylsu/_2742_ ( .A(\mylsu/_0132_ ), .Z(\mylsu/_1264_ ) );
BUF_X1 \mylsu/_2743_ ( .A(\LS_WB_wdata_csreg [1] ), .Z(\mylsu/_0990_ ) );
BUF_X1 \mylsu/_2744_ ( .A(\mylsu/_0133_ ), .Z(\mylsu/_1265_ ) );
BUF_X1 \mylsu/_2745_ ( .A(\LS_WB_wdata_csreg [2] ), .Z(\mylsu/_1001_ ) );
BUF_X1 \mylsu/_2746_ ( .A(\mylsu/_0134_ ), .Z(\mylsu/_1266_ ) );
BUF_X1 \mylsu/_2747_ ( .A(\LS_WB_wdata_csreg [3] ), .Z(\mylsu/_1004_ ) );
BUF_X1 \mylsu/_2748_ ( .A(\mylsu/_0135_ ), .Z(\mylsu/_1267_ ) );
BUF_X1 \mylsu/_2749_ ( .A(\LS_WB_wdata_csreg [4] ), .Z(\mylsu/_1005_ ) );
BUF_X1 \mylsu/_2750_ ( .A(\mylsu/_0136_ ), .Z(\mylsu/_1268_ ) );
BUF_X1 \mylsu/_2751_ ( .A(\LS_WB_wdata_csreg [5] ), .Z(\mylsu/_1006_ ) );
BUF_X1 \mylsu/_2752_ ( .A(\mylsu/_0137_ ), .Z(\mylsu/_1269_ ) );
BUF_X1 \mylsu/_2753_ ( .A(\LS_WB_wdata_csreg [6] ), .Z(\mylsu/_1007_ ) );
BUF_X1 \mylsu/_2754_ ( .A(\mylsu/_0138_ ), .Z(\mylsu/_1270_ ) );
BUF_X1 \mylsu/_2755_ ( .A(\LS_WB_wdata_csreg [7] ), .Z(\mylsu/_1008_ ) );
BUF_X1 \mylsu/_2756_ ( .A(\mylsu/_0139_ ), .Z(\mylsu/_1271_ ) );
BUF_X1 \mylsu/_2757_ ( .A(\LS_WB_wdata_csreg [8] ), .Z(\mylsu/_1009_ ) );
BUF_X1 \mylsu/_2758_ ( .A(\mylsu/_0140_ ), .Z(\mylsu/_1272_ ) );
BUF_X1 \mylsu/_2759_ ( .A(\LS_WB_wdata_csreg [9] ), .Z(\mylsu/_1010_ ) );
BUF_X1 \mylsu/_2760_ ( .A(\mylsu/_0141_ ), .Z(\mylsu/_1273_ ) );
BUF_X1 \mylsu/_2761_ ( .A(\LS_WB_wdata_csreg [10] ), .Z(\mylsu/_0980_ ) );
BUF_X1 \mylsu/_2762_ ( .A(\mylsu/_0142_ ), .Z(\mylsu/_1274_ ) );
BUF_X1 \mylsu/_2763_ ( .A(\LS_WB_wdata_csreg [11] ), .Z(\mylsu/_0981_ ) );
BUF_X1 \mylsu/_2764_ ( .A(\mylsu/_0143_ ), .Z(\mylsu/_1275_ ) );
BUF_X1 \mylsu/_2765_ ( .A(\LS_WB_wdata_csreg [12] ), .Z(\mylsu/_0982_ ) );
BUF_X1 \mylsu/_2766_ ( .A(\mylsu/_0144_ ), .Z(\mylsu/_1276_ ) );
BUF_X1 \mylsu/_2767_ ( .A(\LS_WB_wdata_csreg [13] ), .Z(\mylsu/_0983_ ) );
BUF_X1 \mylsu/_2768_ ( .A(\mylsu/_0145_ ), .Z(\mylsu/_1277_ ) );
BUF_X1 \mylsu/_2769_ ( .A(\LS_WB_wdata_csreg [14] ), .Z(\mylsu/_0984_ ) );
BUF_X1 \mylsu/_2770_ ( .A(\mylsu/_0146_ ), .Z(\mylsu/_1278_ ) );
BUF_X1 \mylsu/_2771_ ( .A(\LS_WB_wdata_csreg [15] ), .Z(\mylsu/_0985_ ) );
BUF_X1 \mylsu/_2772_ ( .A(\mylsu/_0147_ ), .Z(\mylsu/_1279_ ) );
BUF_X1 \mylsu/_2773_ ( .A(\LS_WB_wdata_csreg [16] ), .Z(\mylsu/_0986_ ) );
BUF_X1 \mylsu/_2774_ ( .A(\mylsu/_0148_ ), .Z(\mylsu/_1280_ ) );
BUF_X1 \mylsu/_2775_ ( .A(\LS_WB_wdata_csreg [17] ), .Z(\mylsu/_0987_ ) );
BUF_X1 \mylsu/_2776_ ( .A(\mylsu/_0149_ ), .Z(\mylsu/_1281_ ) );
BUF_X1 \mylsu/_2777_ ( .A(\LS_WB_wdata_csreg [18] ), .Z(\mylsu/_0988_ ) );
BUF_X1 \mylsu/_2778_ ( .A(\mylsu/_0150_ ), .Z(\mylsu/_1282_ ) );
BUF_X1 \mylsu/_2779_ ( .A(\LS_WB_wdata_csreg [19] ), .Z(\mylsu/_0989_ ) );
BUF_X1 \mylsu/_2780_ ( .A(\mylsu/_0151_ ), .Z(\mylsu/_1283_ ) );
BUF_X1 \mylsu/_2781_ ( .A(\LS_WB_wdata_csreg [20] ), .Z(\mylsu/_0991_ ) );
BUF_X1 \mylsu/_2782_ ( .A(\mylsu/_0152_ ), .Z(\mylsu/_1284_ ) );
BUF_X1 \mylsu/_2783_ ( .A(\LS_WB_wdata_csreg [21] ), .Z(\mylsu/_0992_ ) );
BUF_X1 \mylsu/_2784_ ( .A(\mylsu/_0153_ ), .Z(\mylsu/_1285_ ) );
BUF_X1 \mylsu/_2785_ ( .A(\LS_WB_wdata_csreg [22] ), .Z(\mylsu/_0993_ ) );
BUF_X1 \mylsu/_2786_ ( .A(\mylsu/_0154_ ), .Z(\mylsu/_1286_ ) );
BUF_X1 \mylsu/_2787_ ( .A(\LS_WB_wdata_csreg [23] ), .Z(\mylsu/_0994_ ) );
BUF_X1 \mylsu/_2788_ ( .A(\mylsu/_0155_ ), .Z(\mylsu/_1287_ ) );
BUF_X1 \mylsu/_2789_ ( .A(\LS_WB_wdata_csreg [24] ), .Z(\mylsu/_0995_ ) );
BUF_X1 \mylsu/_2790_ ( .A(\mylsu/_0156_ ), .Z(\mylsu/_1288_ ) );
BUF_X1 \mylsu/_2791_ ( .A(\LS_WB_wdata_csreg [25] ), .Z(\mylsu/_0996_ ) );
BUF_X1 \mylsu/_2792_ ( .A(\mylsu/_0157_ ), .Z(\mylsu/_1289_ ) );
BUF_X1 \mylsu/_2793_ ( .A(\LS_WB_wdata_csreg [26] ), .Z(\mylsu/_0997_ ) );
BUF_X1 \mylsu/_2794_ ( .A(\mylsu/_0158_ ), .Z(\mylsu/_1290_ ) );
BUF_X1 \mylsu/_2795_ ( .A(\LS_WB_wdata_csreg [27] ), .Z(\mylsu/_0998_ ) );
BUF_X1 \mylsu/_2796_ ( .A(\mylsu/_0159_ ), .Z(\mylsu/_1291_ ) );
BUF_X1 \mylsu/_2797_ ( .A(\LS_WB_wdata_csreg [28] ), .Z(\mylsu/_0999_ ) );
BUF_X1 \mylsu/_2798_ ( .A(\mylsu/_0160_ ), .Z(\mylsu/_1292_ ) );
BUF_X1 \mylsu/_2799_ ( .A(\LS_WB_wdata_csreg [29] ), .Z(\mylsu/_1000_ ) );
BUF_X1 \mylsu/_2800_ ( .A(\mylsu/_0161_ ), .Z(\mylsu/_1293_ ) );
BUF_X1 \mylsu/_2801_ ( .A(\LS_WB_wdata_csreg [30] ), .Z(\mylsu/_1002_ ) );
BUF_X1 \mylsu/_2802_ ( .A(\mylsu/_0162_ ), .Z(\mylsu/_1294_ ) );
BUF_X1 \mylsu/_2803_ ( .A(\LS_WB_wdata_csreg [31] ), .Z(\mylsu/_1003_ ) );
BUF_X1 \mylsu/_2804_ ( .A(\mylsu/_0163_ ), .Z(\mylsu/_1295_ ) );
BUF_X1 \mylsu/_2805_ ( .A(\mylsu/_0164_ ), .Z(\mylsu/_1296_ ) );
BUF_X1 \mylsu/_2806_ ( .A(\mylsu/_0165_ ), .Z(\mylsu/_1297_ ) );
BUF_X1 \mylsu/_2807_ ( .A(\mylsu/_0166_ ), .Z(\mylsu/_1298_ ) );
BUF_X1 \mylsu/_2808_ ( .A(\mylsu/_0167_ ), .Z(\mylsu/_1299_ ) );
BUF_X1 \mylsu/_2809_ ( .A(\mylsu/_0168_ ), .Z(\mylsu/_1300_ ) );
BUF_X1 \mylsu/_2810_ ( .A(\mylsu/_0169_ ), .Z(\mylsu/_1301_ ) );
BUF_X1 \mylsu/_2811_ ( .A(\mylsu/_0170_ ), .Z(\mylsu/_1302_ ) );
BUF_X1 \mylsu/_2812_ ( .A(\mylsu/_0171_ ), .Z(\mylsu/_1303_ ) );
BUF_X1 \mylsu/_2813_ ( .A(\mylsu/_0172_ ), .Z(\mylsu/_1304_ ) );
BUF_X1 \mylsu/_2814_ ( .A(\mylsu/_0173_ ), .Z(\mylsu/_1305_ ) );
BUF_X1 \mylsu/_2815_ ( .A(\mylsu/_0174_ ), .Z(\mylsu/_1306_ ) );
BUF_X1 \mylsu/_2816_ ( .A(\mylsu/_0175_ ), .Z(\mylsu/_1307_ ) );
BUF_X1 \mylsu/_2817_ ( .A(\mylsu/_0176_ ), .Z(\mylsu/_1308_ ) );
BUF_X1 \mylsu/_2818_ ( .A(\mylsu/_0177_ ), .Z(\mylsu/_1309_ ) );
BUF_X1 \mylsu/_2819_ ( .A(\mylsu/_0178_ ), .Z(\mylsu/_1310_ ) );
BUF_X1 \mylsu/_2820_ ( .A(\mylsu/_0179_ ), .Z(\mylsu/_1311_ ) );
BUF_X1 \mylsu/_2821_ ( .A(\mylsu/_0180_ ), .Z(\mylsu/_1312_ ) );
BUF_X1 \mylsu/_2822_ ( .A(\mylsu/_0181_ ), .Z(\mylsu/_1313_ ) );
BUF_X1 \mylsu/_2823_ ( .A(\mylsu/_0182_ ), .Z(\mylsu/_1314_ ) );
BUF_X1 \mylsu/_2824_ ( .A(\mylsu/_0183_ ), .Z(\mylsu/_1315_ ) );
BUF_X1 \mylsu/_2825_ ( .A(\mylsu/_0184_ ), .Z(\mylsu/_1316_ ) );
BUF_X1 \mylsu/_2826_ ( .A(\mylsu/_0185_ ), .Z(\mylsu/_1317_ ) );
BUF_X1 \mylsu/_2827_ ( .A(\mylsu/_0186_ ), .Z(\mylsu/_1318_ ) );
BUF_X1 \mylsu/_2828_ ( .A(\mylsu/_0187_ ), .Z(\mylsu/_1319_ ) );
BUF_X1 \mylsu/_2829_ ( .A(\mylsu/_0188_ ), .Z(\mylsu/_1320_ ) );
BUF_X1 \mylsu/_2830_ ( .A(\mylsu/_0189_ ), .Z(\mylsu/_1321_ ) );
BUF_X1 \mylsu/_2831_ ( .A(\mylsu/_0190_ ), .Z(\mylsu/_1322_ ) );
BUF_X1 \mylsu/_2832_ ( .A(\mylsu/_0191_ ), .Z(\mylsu/_1323_ ) );
BUF_X1 \mylsu/_2833_ ( .A(\mylsu/_0192_ ), .Z(\mylsu/_1324_ ) );
BUF_X1 \mylsu/_2834_ ( .A(\mylsu/_0193_ ), .Z(\mylsu/_1325_ ) );
BUF_X1 \mylsu/_2835_ ( .A(\mylsu/_0194_ ), .Z(\mylsu/_1326_ ) );
BUF_X1 \mylsu/_2836_ ( .A(\mylsu/_0195_ ), .Z(\mylsu/_1327_ ) );
BUF_X1 \mylsu/_2837_ ( .A(\mylsu/_0196_ ), .Z(\mylsu/_1328_ ) );
BUF_X1 \mylsu/_2838_ ( .A(\mylsu/_0197_ ), .Z(\mylsu/_1329_ ) );
BUF_X1 \mylsu/_2839_ ( .A(\mylsu/_0198_ ), .Z(\mylsu/_1330_ ) );
BUF_X1 \mylsu/_2840_ ( .A(\mylsu/_0199_ ), .Z(\mylsu/_1331_ ) );
BUF_X1 \mylsu/_2841_ ( .A(\mylsu/_0200_ ), .Z(\mylsu/_1332_ ) );
BUF_X1 \mylsu/_2842_ ( .A(\mylsu/_0201_ ), .Z(\mylsu/_1333_ ) );
BUF_X1 \mylsu/_2843_ ( .A(\mylsu/_0202_ ), .Z(\mylsu/_1334_ ) );
BUF_X1 \mylsu/_2844_ ( .A(\mylsu/_0203_ ), .Z(\mylsu/_1335_ ) );
BUF_X1 \mylsu/_2845_ ( .A(\mylsu/_0204_ ), .Z(\mylsu/_1336_ ) );
BUF_X1 \mylsu/_2846_ ( .A(\mylsu/_0205_ ), .Z(\mylsu/_1337_ ) );
BUF_X1 \mylsu/_2847_ ( .A(\mylsu/_0206_ ), .Z(\mylsu/_1338_ ) );
BUF_X1 \mylsu/_2848_ ( .A(\mylsu/_0207_ ), .Z(\mylsu/_1339_ ) );
BUF_X1 \mylsu/_2849_ ( .A(\mylsu/_0208_ ), .Z(\mylsu/_1340_ ) );
BUF_X1 \mylsu/_2850_ ( .A(\mylsu/_0209_ ), .Z(\mylsu/_1341_ ) );
BUF_X1 \mylsu/_2851_ ( .A(\mylsu/_0210_ ), .Z(\mylsu/_1342_ ) );
BUF_X1 \mylsu/_2852_ ( .A(\mylsu/_0211_ ), .Z(\mylsu/_1343_ ) );
BUF_X1 \mylsu/_2853_ ( .A(\mylsu/_0212_ ), .Z(\mylsu/_1344_ ) );
BUF_X1 \mylsu/_2854_ ( .A(\mylsu/_0213_ ), .Z(\mylsu/_1345_ ) );
BUF_X1 \mylsu/_2855_ ( .A(\mylsu/_0214_ ), .Z(\mylsu/_1346_ ) );
BUF_X1 \mylsu/_2856_ ( .A(\mylsu/_0215_ ), .Z(\mylsu/_1347_ ) );
BUF_X1 \mylsu/_2857_ ( .A(\mylsu/_0216_ ), .Z(\mylsu/_1348_ ) );
BUF_X1 \mylsu/_2858_ ( .A(\mylsu/_0217_ ), .Z(\mylsu/_1349_ ) );
BUF_X1 \mylsu/_2859_ ( .A(\mylsu/_0218_ ), .Z(\mylsu/_1350_ ) );
BUF_X1 \mylsu/_2860_ ( .A(\mylsu/_0219_ ), .Z(\mylsu/_1351_ ) );
BUF_X1 \mylsu/_2861_ ( .A(\mylsu/_0220_ ), .Z(\mylsu/_1352_ ) );
BUF_X1 \mylsu/_2862_ ( .A(\mylsu/_0221_ ), .Z(\mylsu/_1353_ ) );
BUF_X1 \mylsu/_2863_ ( .A(\mylsu/_0222_ ), .Z(\mylsu/_1354_ ) );
BUF_X1 \mylsu/_2864_ ( .A(\mylsu/_0223_ ), .Z(\mylsu/_1355_ ) );
BUF_X1 \mylsu/_2865_ ( .A(\mylsu/_0224_ ), .Z(\mylsu/_1356_ ) );
BUF_X1 \mylsu/_2866_ ( .A(\mylsu/_0225_ ), .Z(\mylsu/_1357_ ) );
BUF_X1 \mylsu/_2867_ ( .A(\mylsu/_0226_ ), .Z(\mylsu/_1358_ ) );
BUF_X1 \mylsu/_2868_ ( .A(\mylsu/_0227_ ), .Z(\mylsu/_1359_ ) );
BUF_X1 \mylsu/_2869_ ( .A(\mylsu/_0228_ ), .Z(\mylsu/_1360_ ) );
BUF_X1 \mylsu/_2870_ ( .A(\mylsu/_0229_ ), .Z(\mylsu/_1361_ ) );
BUF_X1 \mylsu/_2871_ ( .A(\mylsu/_0230_ ), .Z(\mylsu/_1362_ ) );
BUF_X1 \mylsu/_2872_ ( .A(\LS_WB_wen_csreg [3] ), .Z(\mylsu/_1043_ ) );
BUF_X1 \mylsu/_2873_ ( .A(\LS_WB_wen_csreg [6] ), .Z(\mylsu/_1044_ ) );
BUF_X1 \mylsu/_2874_ ( .A(\LS_WB_wen_csreg [7] ), .Z(\mylsu/_1045_ ) );
BUF_X1 \mylsu/_2875_ ( .A(\mylsu/_0080_ ), .Z(\mylsu/_1212_ ) );
BUF_X1 \mylsu/_2876_ ( .A(\mylsu/_0130_ ), .Z(\mylsu/_1262_ ) );
BUF_X1 \mylsu/_2877_ ( .A(\mylsu/_0131_ ), .Z(\mylsu/_1263_ ) );
BUF_X1 \mylsu/_2878_ ( .A(\mylsu/_0231_ ), .Z(\mylsu/_1363_ ) );
BUF_X1 \mylsu/_2879_ ( .A(\mylsu/_0232_ ), .Z(\mylsu/_1364_ ) );
BUF_X1 \mylsu/_2880_ ( .A(\mylsu/_0233_ ), .Z(\mylsu/_1365_ ) );
AND2_X1 \myminixbar/_0508_ ( .A1(\myminixbar/_0053_ ), .A2(fanout_net_28 ), .ZN(\myminixbar/_0159_ ) );
NOR2_X4 \myminixbar/_0509_ ( .A1(\myminixbar/_0505_ ), .A2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0160_ ) );
INV_X2 \myminixbar/_0510_ ( .A(\myminixbar/_0485_ ), .ZN(\myminixbar/_0161_ ) );
NOR2_X4 \myminixbar/_0511_ ( .A1(\myminixbar/_0160_ ), .A2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0162_ ) );
MUX2_X1 \myminixbar/_0512_ ( .A(\myminixbar/_0159_ ), .B(\myminixbar/_0021_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0085_ ) );
AND2_X1 \myminixbar/_0513_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0043_ ), .ZN(\myminixbar/_0163_ ) );
MUX2_X1 \myminixbar/_0514_ ( .A(\myminixbar/_0163_ ), .B(\myminixbar/_0011_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0075_ ) );
AND2_X1 \myminixbar/_0515_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0044_ ), .ZN(\myminixbar/_0164_ ) );
MUX2_X1 \myminixbar/_0516_ ( .A(\myminixbar/_0164_ ), .B(\myminixbar/_0012_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0076_ ) );
OAI211_X2 \myminixbar/_0517_ ( .A(fanout_net_28 ), .B(\myminixbar/_0045_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0165_ ) );
OAI211_X2 \myminixbar/_0518_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0013_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0166_ ) );
NAND2_X1 \myminixbar/_0519_ ( .A1(\myminixbar/_0165_ ), .A2(\myminixbar/_0166_ ), .ZN(\myminixbar/_0077_ ) );
OAI211_X2 \myminixbar/_0520_ ( .A(fanout_net_28 ), .B(\myminixbar/_0046_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0167_ ) );
OAI211_X2 \myminixbar/_0521_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0014_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0168_ ) );
NAND2_X1 \myminixbar/_0522_ ( .A1(\myminixbar/_0167_ ), .A2(\myminixbar/_0168_ ), .ZN(\myminixbar/_0078_ ) );
AND2_X1 \myminixbar/_0523_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0048_ ), .ZN(\myminixbar/_0169_ ) );
BUF_X4 \myminixbar/_0524_ ( .A(\myminixbar/_0162_ ), .Z(\myminixbar/_0170_ ) );
MUX2_X1 \myminixbar/_0525_ ( .A(\myminixbar/_0169_ ), .B(\myminixbar/_0016_ ), .S(\myminixbar/_0170_ ), .Z(\myminixbar/_0080_ ) );
AND2_X1 \myminixbar/_0526_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0049_ ), .ZN(\myminixbar/_0171_ ) );
MUX2_X1 \myminixbar/_0527_ ( .A(\myminixbar/_0171_ ), .B(\myminixbar/_0017_ ), .S(\myminixbar/_0170_ ), .Z(\myminixbar/_0081_ ) );
OAI211_X2 \myminixbar/_0528_ ( .A(fanout_net_28 ), .B(\myminixbar/_0050_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0172_ ) );
OAI211_X2 \myminixbar/_0529_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0018_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0173_ ) );
NAND2_X1 \myminixbar/_0530_ ( .A1(\myminixbar/_0172_ ), .A2(\myminixbar/_0173_ ), .ZN(\myminixbar/_0082_ ) );
OAI211_X2 \myminixbar/_0531_ ( .A(fanout_net_28 ), .B(\myminixbar/_0051_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0174_ ) );
OAI211_X2 \myminixbar/_0532_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0019_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0175_ ) );
NAND2_X1 \myminixbar/_0533_ ( .A1(\myminixbar/_0174_ ), .A2(\myminixbar/_0175_ ), .ZN(\myminixbar/_0083_ ) );
OAI211_X2 \myminixbar/_0534_ ( .A(fanout_net_28 ), .B(\myminixbar/_0052_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0176_ ) );
OAI211_X2 \myminixbar/_0535_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0020_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0177_ ) );
NAND2_X1 \myminixbar/_0536_ ( .A1(\myminixbar/_0176_ ), .A2(\myminixbar/_0177_ ), .ZN(\myminixbar/_0084_ ) );
AND2_X1 \myminixbar/_0537_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0054_ ), .ZN(\myminixbar/_0178_ ) );
MUX2_X1 \myminixbar/_0538_ ( .A(\myminixbar/_0178_ ), .B(\myminixbar/_0022_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0086_ ) );
AND2_X1 \myminixbar/_0539_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0055_ ), .ZN(\myminixbar/_0179_ ) );
MUX2_X1 \myminixbar/_0540_ ( .A(\myminixbar/_0179_ ), .B(\myminixbar/_0023_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0087_ ) );
AND2_X1 \myminixbar/_0541_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0056_ ), .ZN(\myminixbar/_0180_ ) );
MUX2_X1 \myminixbar/_0542_ ( .A(\myminixbar/_0180_ ), .B(\myminixbar/_0024_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0088_ ) );
AND2_X1 \myminixbar/_0543_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0057_ ), .ZN(\myminixbar/_0181_ ) );
MUX2_X1 \myminixbar/_0544_ ( .A(\myminixbar/_0181_ ), .B(\myminixbar/_0025_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0089_ ) );
AND2_X1 \myminixbar/_0545_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0059_ ), .ZN(\myminixbar/_0182_ ) );
MUX2_X1 \myminixbar/_0546_ ( .A(\myminixbar/_0182_ ), .B(\myminixbar/_0027_ ), .S(\myminixbar/_0170_ ), .Z(\myminixbar/_0091_ ) );
AND2_X1 \myminixbar/_0547_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0060_ ), .ZN(\myminixbar/_0183_ ) );
MUX2_X1 \myminixbar/_0548_ ( .A(\myminixbar/_0183_ ), .B(\myminixbar/_0028_ ), .S(\myminixbar/_0162_ ), .Z(\myminixbar/_0092_ ) );
NAND4_X1 \myminixbar/_0549_ ( .A1(\myminixbar/_0174_ ), .A2(\myminixbar/_0176_ ), .A3(\myminixbar/_0175_ ), .A4(\myminixbar/_0177_ ), .ZN(\myminixbar/_0184_ ) );
OR3_X1 \myminixbar/_0550_ ( .A1(\myminixbar/_0086_ ), .A2(\myminixbar/_0087_ ), .A3(\myminixbar/_0184_ ), .ZN(\myminixbar/_0185_ ) );
OR2_X1 \myminixbar/_0551_ ( .A1(\myminixbar/_0088_ ), .A2(\myminixbar/_0089_ ), .ZN(\myminixbar/_0186_ ) );
OR4_X4 \myminixbar/_0552_ ( .A1(\myminixbar/_0091_ ), .A2(\myminixbar/_0185_ ), .A3(\myminixbar/_0092_ ), .A4(\myminixbar/_0186_ ), .ZN(\myminixbar/_0187_ ) );
NAND3_X1 \myminixbar/_0553_ ( .A1(\myminixbar/_0085_ ), .A2(\myminixbar/_0165_ ), .A3(\myminixbar/_0166_ ), .ZN(\myminixbar/_0188_ ) );
OR3_X1 \myminixbar/_0554_ ( .A1(\myminixbar/_0188_ ), .A2(\myminixbar/_0075_ ), .A3(\myminixbar/_0076_ ), .ZN(\myminixbar/_0189_ ) );
NAND4_X1 \myminixbar/_0555_ ( .A1(\myminixbar/_0167_ ), .A2(\myminixbar/_0172_ ), .A3(\myminixbar/_0168_ ), .A4(\myminixbar/_0173_ ), .ZN(\myminixbar/_0190_ ) );
OR4_X4 \myminixbar/_0556_ ( .A1(\myminixbar/_0080_ ), .A2(\myminixbar/_0189_ ), .A3(\myminixbar/_0081_ ), .A4(\myminixbar/_0190_ ), .ZN(\myminixbar/_0191_ ) );
OAI211_X2 \myminixbar/_0557_ ( .A(fanout_net_28 ), .B(\myminixbar/_0156_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0192_ ) );
OAI211_X2 \myminixbar/_0558_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0155_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0193_ ) );
AND2_X1 \myminixbar/_0559_ ( .A1(\myminixbar/_0192_ ), .A2(\myminixbar/_0193_ ), .ZN(\myminixbar/_0194_ ) );
NOR3_X1 \myminixbar/_0560_ ( .A1(\myminixbar/_0187_ ), .A2(\myminixbar/_0191_ ), .A3(\myminixbar/_0194_ ), .ZN(\myminixbar/_0157_ ) );
OR3_X1 \myminixbar/_0561_ ( .A1(\myminixbar/_0191_ ), .A2(\myminixbar/_0144_ ), .A3(\myminixbar/_0187_ ), .ZN(\myminixbar/_0195_ ) );
NOR2_X4 \myminixbar/_0562_ ( .A1(\myminixbar/_0191_ ), .A2(\myminixbar/_0187_ ), .ZN(\myminixbar/_0196_ ) );
BUF_X4 \myminixbar/_0563_ ( .A(\myminixbar/_0196_ ), .Z(\myminixbar/_0197_ ) );
OAI21_X1 \myminixbar/_0564_ ( .A(\myminixbar/_0195_ ), .B1(\myminixbar/_0145_ ), .B2(\myminixbar/_0197_ ), .ZN(\myminixbar/_0198_ ) );
INV_X2 \myminixbar/_0565_ ( .A(\myminixbar/_0170_ ), .ZN(\myminixbar/_0199_ ) );
BUF_X4 \myminixbar/_0566_ ( .A(\myminixbar/_0199_ ), .Z(\myminixbar/_0200_ ) );
NOR2_X1 \myminixbar/_0567_ ( .A1(\myminixbar/_0198_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0142_ ) );
NAND2_X2 \myminixbar/_0568_ ( .A1(\myminixbar/_0199_ ), .A2(fanout_net_28 ), .ZN(\myminixbar/_0201_ ) );
BUF_X4 \myminixbar/_0569_ ( .A(\myminixbar/_0201_ ), .Z(\myminixbar/_0202_ ) );
NOR2_X1 \myminixbar/_0570_ ( .A1(\myminixbar/_0198_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0143_ ) );
AND2_X4 \myminixbar/_0571_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0502_ ), .ZN(\myminixbar/_0203_ ) );
INV_X4 \myminixbar/_0572_ ( .A(\myminixbar/_0196_ ), .ZN(\myminixbar/_0204_ ) );
BUF_X4 \myminixbar/_0573_ ( .A(\myminixbar/_0204_ ), .Z(\myminixbar/_0205_ ) );
AOI21_X2 \myminixbar/_0574_ ( .A(\myminixbar/_0203_ ), .B1(\myminixbar/_0503_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0206_ ) );
NOR2_X1 \myminixbar/_0575_ ( .A1(\myminixbar/_0206_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0500_ ) );
NOR2_X1 \myminixbar/_0576_ ( .A1(\myminixbar/_0206_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0501_ ) );
OAI211_X2 \myminixbar/_0577_ ( .A(fanout_net_28 ), .B(\myminixbar/_0488_ ), .C1(\myminixbar/_0160_ ), .C2(\myminixbar/_0161_ ), .ZN(\myminixbar/_0207_ ) );
OAI211_X2 \myminixbar/_0578_ ( .A(\myminixbar/_0485_ ), .B(\myminixbar/_0487_ ), .C1(\myminixbar/_0505_ ), .C2(\myminixbar/_0504_ ), .ZN(\myminixbar/_0208_ ) );
AND2_X1 \myminixbar/_0579_ ( .A1(\myminixbar/_0207_ ), .A2(\myminixbar/_0208_ ), .ZN(\myminixbar/_0209_ ) );
NOR3_X1 \myminixbar/_0580_ ( .A1(\myminixbar/_0187_ ), .A2(\myminixbar/_0191_ ), .A3(\myminixbar/_0209_ ), .ZN(\myminixbar/_0489_ ) );
AND2_X4 \myminixbar/_0581_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0483_ ), .ZN(\myminixbar/_0210_ ) );
AOI21_X2 \myminixbar/_0582_ ( .A(\myminixbar/_0210_ ), .B1(\myminixbar/_0484_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0211_ ) );
NOR2_X1 \myminixbar/_0583_ ( .A1(\myminixbar/_0211_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0481_ ) );
NOR2_X1 \myminixbar/_0584_ ( .A1(\myminixbar/_0211_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0482_ ) );
INV_X1 \myminixbar/_0585_ ( .A(\myminixbar/_0499_ ), .ZN(\myminixbar/_0212_ ) );
OAI21_X1 \myminixbar/_0586_ ( .A(\myminixbar/_0212_ ), .B1(fanout_net_28 ), .B2(\myminixbar/_0485_ ), .ZN(\myminixbar/_0002_ ) );
AOI211_X4 \myminixbar/_0587_ ( .A(\myminixbar/_0499_ ), .B(\myminixbar/_0161_ ), .C1(\myminixbar/_0160_ ), .C2(fanout_net_28 ), .ZN(\myminixbar/_0003_ ) );
AND2_X1 \myminixbar/_0588_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0036_ ), .ZN(\myminixbar/_0213_ ) );
BUF_X4 \myminixbar/_0589_ ( .A(\myminixbar/_0170_ ), .Z(\myminixbar/_0214_ ) );
MUX2_X1 \myminixbar/_0590_ ( .A(\myminixbar/_0213_ ), .B(\myminixbar/_0004_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0068_ ) );
AND2_X1 \myminixbar/_0591_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0047_ ), .ZN(\myminixbar/_0215_ ) );
MUX2_X1 \myminixbar/_0592_ ( .A(\myminixbar/_0215_ ), .B(\myminixbar/_0015_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0079_ ) );
AND2_X1 \myminixbar/_0593_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0058_ ), .ZN(\myminixbar/_0216_ ) );
MUX2_X1 \myminixbar/_0594_ ( .A(\myminixbar/_0216_ ), .B(\myminixbar/_0026_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0090_ ) );
AND2_X1 \myminixbar/_0595_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0061_ ), .ZN(\myminixbar/_0217_ ) );
MUX2_X1 \myminixbar/_0596_ ( .A(\myminixbar/_0217_ ), .B(\myminixbar/_0029_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0093_ ) );
AND2_X1 \myminixbar/_0597_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0062_ ), .ZN(\myminixbar/_0218_ ) );
MUX2_X1 \myminixbar/_0598_ ( .A(\myminixbar/_0218_ ), .B(\myminixbar/_0030_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0094_ ) );
AND2_X1 \myminixbar/_0599_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0063_ ), .ZN(\myminixbar/_0219_ ) );
MUX2_X1 \myminixbar/_0600_ ( .A(\myminixbar/_0219_ ), .B(\myminixbar/_0031_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0095_ ) );
AND2_X1 \myminixbar/_0601_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0064_ ), .ZN(\myminixbar/_0220_ ) );
MUX2_X1 \myminixbar/_0602_ ( .A(\myminixbar/_0220_ ), .B(\myminixbar/_0032_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0096_ ) );
AND2_X1 \myminixbar/_0603_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0065_ ), .ZN(\myminixbar/_0221_ ) );
MUX2_X1 \myminixbar/_0604_ ( .A(\myminixbar/_0221_ ), .B(\myminixbar/_0033_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0097_ ) );
AND2_X1 \myminixbar/_0605_ ( .A1(fanout_net_28 ), .A2(\myminixbar/_0066_ ), .ZN(\myminixbar/_0222_ ) );
MUX2_X1 \myminixbar/_0606_ ( .A(\myminixbar/_0222_ ), .B(\myminixbar/_0034_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0098_ ) );
AND2_X1 \myminixbar/_0607_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0067_ ), .ZN(\myminixbar/_0223_ ) );
MUX2_X1 \myminixbar/_0608_ ( .A(\myminixbar/_0223_ ), .B(\myminixbar/_0035_ ), .S(\myminixbar/_0214_ ), .Z(\myminixbar/_0099_ ) );
AND2_X1 \myminixbar/_0609_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0037_ ), .ZN(\myminixbar/_0224_ ) );
BUF_X4 \myminixbar/_0610_ ( .A(\myminixbar/_0170_ ), .Z(\myminixbar/_0225_ ) );
MUX2_X1 \myminixbar/_0611_ ( .A(\myminixbar/_0224_ ), .B(\myminixbar/_0005_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0069_ ) );
AND2_X1 \myminixbar/_0612_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0038_ ), .ZN(\myminixbar/_0226_ ) );
MUX2_X1 \myminixbar/_0613_ ( .A(\myminixbar/_0226_ ), .B(\myminixbar/_0006_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0070_ ) );
AND2_X1 \myminixbar/_0614_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0039_ ), .ZN(\myminixbar/_0227_ ) );
MUX2_X1 \myminixbar/_0615_ ( .A(\myminixbar/_0227_ ), .B(\myminixbar/_0007_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0071_ ) );
AND2_X1 \myminixbar/_0616_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0040_ ), .ZN(\myminixbar/_0228_ ) );
MUX2_X1 \myminixbar/_0617_ ( .A(\myminixbar/_0228_ ), .B(\myminixbar/_0008_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0072_ ) );
AND2_X1 \myminixbar/_0618_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0041_ ), .ZN(\myminixbar/_0229_ ) );
MUX2_X1 \myminixbar/_0619_ ( .A(\myminixbar/_0229_ ), .B(\myminixbar/_0009_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0073_ ) );
AND2_X1 \myminixbar/_0620_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0042_ ), .ZN(\myminixbar/_0230_ ) );
MUX2_X1 \myminixbar/_0621_ ( .A(\myminixbar/_0230_ ), .B(\myminixbar/_0010_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0074_ ) );
NOR2_X1 \myminixbar/_0622_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0194_ ), .ZN(\myminixbar/_0158_ ) );
AND2_X1 \myminixbar/_0623_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0110_ ), .ZN(\myminixbar/_0231_ ) );
MUX2_X1 \myminixbar/_0624_ ( .A(\myminixbar/_0231_ ), .B(\myminixbar/_0106_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0114_ ) );
AND2_X1 \myminixbar/_0625_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0111_ ), .ZN(\myminixbar/_0232_ ) );
MUX2_X1 \myminixbar/_0626_ ( .A(\myminixbar/_0232_ ), .B(\myminixbar/_0107_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0115_ ) );
AND2_X1 \myminixbar/_0627_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0112_ ), .ZN(\myminixbar/_0233_ ) );
MUX2_X1 \myminixbar/_0628_ ( .A(\myminixbar/_0233_ ), .B(\myminixbar/_0108_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0116_ ) );
AND2_X1 \myminixbar/_0629_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0113_ ), .ZN(\myminixbar/_0234_ ) );
MUX2_X1 \myminixbar/_0630_ ( .A(\myminixbar/_0234_ ), .B(\myminixbar/_0109_ ), .S(\myminixbar/_0225_ ), .Z(\myminixbar/_0117_ ) );
AND2_X1 \myminixbar/_0631_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0126_ ), .ZN(\myminixbar/_0235_ ) );
BUF_X4 \myminixbar/_0632_ ( .A(\myminixbar/_0170_ ), .Z(\myminixbar/_0236_ ) );
MUX2_X1 \myminixbar/_0633_ ( .A(\myminixbar/_0235_ ), .B(\myminixbar/_0118_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0134_ ) );
AND2_X1 \myminixbar/_0634_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0127_ ), .ZN(\myminixbar/_0237_ ) );
MUX2_X1 \myminixbar/_0635_ ( .A(\myminixbar/_0237_ ), .B(\myminixbar/_0119_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0135_ ) );
AND2_X1 \myminixbar/_0636_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0128_ ), .ZN(\myminixbar/_0238_ ) );
MUX2_X1 \myminixbar/_0637_ ( .A(\myminixbar/_0238_ ), .B(\myminixbar/_0120_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0136_ ) );
AND2_X1 \myminixbar/_0638_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0129_ ), .ZN(\myminixbar/_0239_ ) );
MUX2_X1 \myminixbar/_0639_ ( .A(\myminixbar/_0239_ ), .B(\myminixbar/_0121_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0137_ ) );
AND2_X1 \myminixbar/_0640_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0130_ ), .ZN(\myminixbar/_0240_ ) );
MUX2_X1 \myminixbar/_0641_ ( .A(\myminixbar/_0240_ ), .B(\myminixbar/_0122_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0138_ ) );
AND2_X1 \myminixbar/_0642_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0131_ ), .ZN(\myminixbar/_0241_ ) );
MUX2_X1 \myminixbar/_0643_ ( .A(\myminixbar/_0241_ ), .B(\myminixbar/_0123_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0139_ ) );
AND2_X1 \myminixbar/_0644_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0132_ ), .ZN(\myminixbar/_0242_ ) );
MUX2_X1 \myminixbar/_0645_ ( .A(\myminixbar/_0242_ ), .B(\myminixbar/_0124_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0140_ ) );
AND2_X1 \myminixbar/_0646_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0133_ ), .ZN(\myminixbar/_0243_ ) );
MUX2_X1 \myminixbar/_0647_ ( .A(\myminixbar/_0243_ ), .B(\myminixbar/_0125_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0141_ ) );
AND2_X1 \myminixbar/_0648_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0149_ ), .ZN(\myminixbar/_0244_ ) );
MUX2_X1 \myminixbar/_0649_ ( .A(\myminixbar/_0244_ ), .B(\myminixbar/_0146_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0152_ ) );
AND2_X1 \myminixbar/_0650_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0150_ ), .ZN(\myminixbar/_0245_ ) );
MUX2_X1 \myminixbar/_0651_ ( .A(\myminixbar/_0245_ ), .B(\myminixbar/_0147_ ), .S(\myminixbar/_0236_ ), .Z(\myminixbar/_0153_ ) );
AND2_X1 \myminixbar/_0652_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0151_ ), .ZN(\myminixbar/_0246_ ) );
MUX2_X1 \myminixbar/_0653_ ( .A(\myminixbar/_0246_ ), .B(\myminixbar/_0148_ ), .S(\myminixbar/_0170_ ), .Z(\myminixbar/_0154_ ) );
AND2_X1 \myminixbar/_0654_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0102_ ), .ZN(\myminixbar/_0247_ ) );
MUX2_X1 \myminixbar/_0655_ ( .A(\myminixbar/_0247_ ), .B(\myminixbar/_0100_ ), .S(\myminixbar/_0170_ ), .Z(\myminixbar/_0104_ ) );
AND2_X1 \myminixbar/_0656_ ( .A1(\myminixbar/_0486_ ), .A2(\myminixbar/_0103_ ), .ZN(\myminixbar/_0248_ ) );
MUX2_X1 \myminixbar/_0657_ ( .A(\myminixbar/_0248_ ), .B(\myminixbar/_0101_ ), .S(\myminixbar/_0170_ ), .Z(\myminixbar/_0105_ ) );
AND2_X4 \myminixbar/_0658_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0401_ ), .ZN(\myminixbar/_0249_ ) );
AOI21_X2 \myminixbar/_0659_ ( .A(\myminixbar/_0249_ ), .B1(\myminixbar/_0433_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0250_ ) );
NOR2_X1 \myminixbar/_0660_ ( .A1(\myminixbar/_0250_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0337_ ) );
AND2_X4 \myminixbar/_0661_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0412_ ), .ZN(\myminixbar/_0251_ ) );
AOI21_X2 \myminixbar/_0662_ ( .A(\myminixbar/_0251_ ), .B1(\myminixbar/_0444_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0252_ ) );
NOR2_X1 \myminixbar/_0663_ ( .A1(\myminixbar/_0252_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0348_ ) );
AND2_X4 \myminixbar/_0664_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0423_ ), .ZN(\myminixbar/_0253_ ) );
AOI21_X2 \myminixbar/_0665_ ( .A(\myminixbar/_0253_ ), .B1(\myminixbar/_0455_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0254_ ) );
NOR2_X1 \myminixbar/_0666_ ( .A1(\myminixbar/_0254_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0359_ ) );
AND2_X4 \myminixbar/_0667_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0426_ ), .ZN(\myminixbar/_0255_ ) );
AOI21_X2 \myminixbar/_0668_ ( .A(\myminixbar/_0255_ ), .B1(\myminixbar/_0458_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0256_ ) );
NOR2_X1 \myminixbar/_0669_ ( .A1(\myminixbar/_0256_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0362_ ) );
AND2_X4 \myminixbar/_0670_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0427_ ), .ZN(\myminixbar/_0257_ ) );
AOI21_X2 \myminixbar/_0671_ ( .A(\myminixbar/_0257_ ), .B1(\myminixbar/_0459_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0258_ ) );
NOR2_X1 \myminixbar/_0672_ ( .A1(\myminixbar/_0258_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0363_ ) );
BUF_X4 \myminixbar/_0673_ ( .A(\myminixbar/_0196_ ), .Z(\myminixbar/_0259_ ) );
AND2_X1 \myminixbar/_0674_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0428_ ), .ZN(\myminixbar/_0260_ ) );
AOI21_X1 \myminixbar/_0675_ ( .A(\myminixbar/_0260_ ), .B1(\myminixbar/_0460_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0261_ ) );
NOR2_X1 \myminixbar/_0676_ ( .A1(\myminixbar/_0261_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0364_ ) );
AND2_X1 \myminixbar/_0677_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0429_ ), .ZN(\myminixbar/_0262_ ) );
AOI21_X1 \myminixbar/_0678_ ( .A(\myminixbar/_0262_ ), .B1(\myminixbar/_0461_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0263_ ) );
NOR2_X1 \myminixbar/_0679_ ( .A1(\myminixbar/_0263_ ), .A2(\myminixbar/_0200_ ), .ZN(\myminixbar/_0365_ ) );
AND2_X1 \myminixbar/_0680_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0430_ ), .ZN(\myminixbar/_0264_ ) );
AOI21_X1 \myminixbar/_0681_ ( .A(\myminixbar/_0264_ ), .B1(\myminixbar/_0462_ ), .B2(\myminixbar/_0205_ ), .ZN(\myminixbar/_0265_ ) );
BUF_X4 \myminixbar/_0682_ ( .A(\myminixbar/_0199_ ), .Z(\myminixbar/_0266_ ) );
NOR2_X1 \myminixbar/_0683_ ( .A1(\myminixbar/_0265_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0366_ ) );
AND2_X1 \myminixbar/_0684_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0431_ ), .ZN(\myminixbar/_0267_ ) );
BUF_X4 \myminixbar/_0685_ ( .A(\myminixbar/_0204_ ), .Z(\myminixbar/_0268_ ) );
AOI21_X2 \myminixbar/_0686_ ( .A(\myminixbar/_0267_ ), .B1(\myminixbar/_0463_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0269_ ) );
NOR2_X1 \myminixbar/_0687_ ( .A1(\myminixbar/_0269_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0367_ ) );
AND2_X1 \myminixbar/_0688_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0432_ ), .ZN(\myminixbar/_0270_ ) );
AOI21_X2 \myminixbar/_0689_ ( .A(\myminixbar/_0270_ ), .B1(\myminixbar/_0464_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0271_ ) );
NOR2_X1 \myminixbar/_0690_ ( .A1(\myminixbar/_0271_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0368_ ) );
AND2_X1 \myminixbar/_0691_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0402_ ), .ZN(\myminixbar/_0272_ ) );
AOI21_X2 \myminixbar/_0692_ ( .A(\myminixbar/_0272_ ), .B1(\myminixbar/_0434_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0273_ ) );
NOR2_X1 \myminixbar/_0693_ ( .A1(\myminixbar/_0273_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0338_ ) );
AND2_X1 \myminixbar/_0694_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0403_ ), .ZN(\myminixbar/_0274_ ) );
AOI21_X2 \myminixbar/_0695_ ( .A(\myminixbar/_0274_ ), .B1(\myminixbar/_0435_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0275_ ) );
NOR2_X1 \myminixbar/_0696_ ( .A1(\myminixbar/_0275_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0339_ ) );
AND2_X1 \myminixbar/_0697_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0404_ ), .ZN(\myminixbar/_0276_ ) );
AOI21_X2 \myminixbar/_0698_ ( .A(\myminixbar/_0276_ ), .B1(\myminixbar/_0436_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0277_ ) );
NOR2_X1 \myminixbar/_0699_ ( .A1(\myminixbar/_0277_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0340_ ) );
AND2_X1 \myminixbar/_0700_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0405_ ), .ZN(\myminixbar/_0278_ ) );
AOI21_X2 \myminixbar/_0701_ ( .A(\myminixbar/_0278_ ), .B1(\myminixbar/_0437_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0279_ ) );
NOR2_X1 \myminixbar/_0702_ ( .A1(\myminixbar/_0279_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0341_ ) );
AND2_X1 \myminixbar/_0703_ ( .A1(\myminixbar/_0259_ ), .A2(\myminixbar/_0406_ ), .ZN(\myminixbar/_0280_ ) );
AOI21_X2 \myminixbar/_0704_ ( .A(\myminixbar/_0280_ ), .B1(\myminixbar/_0438_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0281_ ) );
NOR2_X1 \myminixbar/_0705_ ( .A1(\myminixbar/_0281_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0342_ ) );
BUF_X4 \myminixbar/_0706_ ( .A(\myminixbar/_0196_ ), .Z(\myminixbar/_0282_ ) );
AND2_X1 \myminixbar/_0707_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0407_ ), .ZN(\myminixbar/_0283_ ) );
AOI21_X2 \myminixbar/_0708_ ( .A(\myminixbar/_0283_ ), .B1(\myminixbar/_0439_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0284_ ) );
NOR2_X1 \myminixbar/_0709_ ( .A1(\myminixbar/_0284_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0343_ ) );
AND2_X1 \myminixbar/_0710_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0408_ ), .ZN(\myminixbar/_0285_ ) );
AOI21_X2 \myminixbar/_0711_ ( .A(\myminixbar/_0285_ ), .B1(\myminixbar/_0440_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0286_ ) );
NOR2_X1 \myminixbar/_0712_ ( .A1(\myminixbar/_0286_ ), .A2(\myminixbar/_0266_ ), .ZN(\myminixbar/_0344_ ) );
AND2_X1 \myminixbar/_0713_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0409_ ), .ZN(\myminixbar/_0287_ ) );
AOI21_X2 \myminixbar/_0714_ ( .A(\myminixbar/_0287_ ), .B1(\myminixbar/_0441_ ), .B2(\myminixbar/_0268_ ), .ZN(\myminixbar/_0288_ ) );
BUF_X4 \myminixbar/_0715_ ( .A(\myminixbar/_0199_ ), .Z(\myminixbar/_0289_ ) );
NOR2_X1 \myminixbar/_0716_ ( .A1(\myminixbar/_0288_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0345_ ) );
AND2_X1 \myminixbar/_0717_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0410_ ), .ZN(\myminixbar/_0290_ ) );
BUF_X4 \myminixbar/_0718_ ( .A(\myminixbar/_0204_ ), .Z(\myminixbar/_0291_ ) );
AOI21_X1 \myminixbar/_0719_ ( .A(\myminixbar/_0290_ ), .B1(\myminixbar/_0442_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0292_ ) );
NOR2_X1 \myminixbar/_0720_ ( .A1(\myminixbar/_0292_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0346_ ) );
AND2_X1 \myminixbar/_0721_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0411_ ), .ZN(\myminixbar/_0293_ ) );
AOI21_X1 \myminixbar/_0722_ ( .A(\myminixbar/_0293_ ), .B1(\myminixbar/_0443_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0294_ ) );
NOR2_X1 \myminixbar/_0723_ ( .A1(\myminixbar/_0294_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0347_ ) );
AND2_X1 \myminixbar/_0724_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0413_ ), .ZN(\myminixbar/_0295_ ) );
AOI21_X1 \myminixbar/_0725_ ( .A(\myminixbar/_0295_ ), .B1(\myminixbar/_0445_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0296_ ) );
NOR2_X1 \myminixbar/_0726_ ( .A1(\myminixbar/_0296_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0349_ ) );
AND2_X1 \myminixbar/_0727_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0414_ ), .ZN(\myminixbar/_0297_ ) );
AOI21_X2 \myminixbar/_0728_ ( .A(\myminixbar/_0297_ ), .B1(\myminixbar/_0446_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0298_ ) );
NOR2_X1 \myminixbar/_0729_ ( .A1(\myminixbar/_0298_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0350_ ) );
AND2_X1 \myminixbar/_0730_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0415_ ), .ZN(\myminixbar/_0299_ ) );
AOI21_X1 \myminixbar/_0731_ ( .A(\myminixbar/_0299_ ), .B1(\myminixbar/_0447_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0300_ ) );
NOR2_X1 \myminixbar/_0732_ ( .A1(\myminixbar/_0300_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0351_ ) );
AND2_X1 \myminixbar/_0733_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0416_ ), .ZN(\myminixbar/_0301_ ) );
AOI21_X1 \myminixbar/_0734_ ( .A(\myminixbar/_0301_ ), .B1(\myminixbar/_0448_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0302_ ) );
NOR2_X1 \myminixbar/_0735_ ( .A1(\myminixbar/_0302_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0352_ ) );
AND2_X1 \myminixbar/_0736_ ( .A1(\myminixbar/_0282_ ), .A2(\myminixbar/_0417_ ), .ZN(\myminixbar/_0303_ ) );
AOI21_X2 \myminixbar/_0737_ ( .A(\myminixbar/_0303_ ), .B1(\myminixbar/_0449_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0304_ ) );
NOR2_X1 \myminixbar/_0738_ ( .A1(\myminixbar/_0304_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0353_ ) );
BUF_X4 \myminixbar/_0739_ ( .A(\myminixbar/_0196_ ), .Z(\myminixbar/_0305_ ) );
AND2_X1 \myminixbar/_0740_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0418_ ), .ZN(\myminixbar/_0306_ ) );
AOI21_X2 \myminixbar/_0741_ ( .A(\myminixbar/_0306_ ), .B1(\myminixbar/_0450_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0307_ ) );
NOR2_X1 \myminixbar/_0742_ ( .A1(\myminixbar/_0307_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0354_ ) );
AND2_X1 \myminixbar/_0743_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0419_ ), .ZN(\myminixbar/_0308_ ) );
AOI21_X2 \myminixbar/_0744_ ( .A(\myminixbar/_0308_ ), .B1(\myminixbar/_0451_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0309_ ) );
NOR2_X1 \myminixbar/_0745_ ( .A1(\myminixbar/_0309_ ), .A2(\myminixbar/_0289_ ), .ZN(\myminixbar/_0355_ ) );
AND2_X1 \myminixbar/_0746_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0420_ ), .ZN(\myminixbar/_0310_ ) );
AOI21_X2 \myminixbar/_0747_ ( .A(\myminixbar/_0310_ ), .B1(\myminixbar/_0452_ ), .B2(\myminixbar/_0291_ ), .ZN(\myminixbar/_0311_ ) );
BUF_X4 \myminixbar/_0748_ ( .A(\myminixbar/_0199_ ), .Z(\myminixbar/_0312_ ) );
NOR2_X1 \myminixbar/_0749_ ( .A1(\myminixbar/_0311_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0356_ ) );
AND2_X1 \myminixbar/_0750_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0421_ ), .ZN(\myminixbar/_0313_ ) );
BUF_X4 \myminixbar/_0751_ ( .A(\myminixbar/_0204_ ), .Z(\myminixbar/_0314_ ) );
AOI21_X2 \myminixbar/_0752_ ( .A(\myminixbar/_0313_ ), .B1(\myminixbar/_0453_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0315_ ) );
NOR2_X1 \myminixbar/_0753_ ( .A1(\myminixbar/_0315_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0357_ ) );
AND2_X1 \myminixbar/_0754_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0422_ ), .ZN(\myminixbar/_0316_ ) );
AOI21_X2 \myminixbar/_0755_ ( .A(\myminixbar/_0316_ ), .B1(\myminixbar/_0454_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0317_ ) );
NOR2_X1 \myminixbar/_0756_ ( .A1(\myminixbar/_0317_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0358_ ) );
AND2_X1 \myminixbar/_0757_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0424_ ), .ZN(\myminixbar/_0318_ ) );
AOI21_X2 \myminixbar/_0758_ ( .A(\myminixbar/_0318_ ), .B1(\myminixbar/_0456_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0319_ ) );
NOR2_X1 \myminixbar/_0759_ ( .A1(\myminixbar/_0319_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0360_ ) );
AND2_X1 \myminixbar/_0760_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0425_ ), .ZN(\myminixbar/_0320_ ) );
AOI21_X2 \myminixbar/_0761_ ( .A(\myminixbar/_0320_ ), .B1(\myminixbar/_0457_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0321_ ) );
NOR2_X1 \myminixbar/_0762_ ( .A1(\myminixbar/_0321_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0361_ ) );
NOR2_X1 \myminixbar/_0763_ ( .A1(\myminixbar/_0250_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0369_ ) );
NOR2_X1 \myminixbar/_0764_ ( .A1(\myminixbar/_0252_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0380_ ) );
NOR2_X1 \myminixbar/_0765_ ( .A1(\myminixbar/_0254_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0391_ ) );
NOR2_X1 \myminixbar/_0766_ ( .A1(\myminixbar/_0256_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0394_ ) );
NOR2_X1 \myminixbar/_0767_ ( .A1(\myminixbar/_0258_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0395_ ) );
NOR2_X1 \myminixbar/_0768_ ( .A1(\myminixbar/_0261_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0396_ ) );
NOR2_X1 \myminixbar/_0769_ ( .A1(\myminixbar/_0263_ ), .A2(\myminixbar/_0202_ ), .ZN(\myminixbar/_0397_ ) );
BUF_X4 \myminixbar/_0770_ ( .A(\myminixbar/_0201_ ), .Z(\myminixbar/_0322_ ) );
NOR2_X1 \myminixbar/_0771_ ( .A1(\myminixbar/_0265_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0398_ ) );
NOR2_X1 \myminixbar/_0772_ ( .A1(\myminixbar/_0269_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0399_ ) );
NOR2_X1 \myminixbar/_0773_ ( .A1(\myminixbar/_0271_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0400_ ) );
NOR2_X1 \myminixbar/_0774_ ( .A1(\myminixbar/_0273_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0370_ ) );
NOR2_X1 \myminixbar/_0775_ ( .A1(\myminixbar/_0275_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0371_ ) );
NOR2_X1 \myminixbar/_0776_ ( .A1(\myminixbar/_0277_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0372_ ) );
NOR2_X1 \myminixbar/_0777_ ( .A1(\myminixbar/_0279_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0373_ ) );
NOR2_X1 \myminixbar/_0778_ ( .A1(\myminixbar/_0281_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0374_ ) );
NOR2_X1 \myminixbar/_0779_ ( .A1(\myminixbar/_0284_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0375_ ) );
NOR2_X1 \myminixbar/_0780_ ( .A1(\myminixbar/_0286_ ), .A2(\myminixbar/_0322_ ), .ZN(\myminixbar/_0376_ ) );
BUF_X4 \myminixbar/_0781_ ( .A(\myminixbar/_0201_ ), .Z(\myminixbar/_0323_ ) );
NOR2_X1 \myminixbar/_0782_ ( .A1(\myminixbar/_0288_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0377_ ) );
NOR2_X1 \myminixbar/_0783_ ( .A1(\myminixbar/_0292_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0378_ ) );
NOR2_X1 \myminixbar/_0784_ ( .A1(\myminixbar/_0294_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0379_ ) );
NOR2_X1 \myminixbar/_0785_ ( .A1(\myminixbar/_0296_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0381_ ) );
NOR2_X1 \myminixbar/_0786_ ( .A1(\myminixbar/_0298_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0382_ ) );
NOR2_X1 \myminixbar/_0787_ ( .A1(\myminixbar/_0300_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0383_ ) );
NOR2_X1 \myminixbar/_0788_ ( .A1(\myminixbar/_0302_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0384_ ) );
NOR2_X1 \myminixbar/_0789_ ( .A1(\myminixbar/_0304_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0385_ ) );
NOR2_X1 \myminixbar/_0790_ ( .A1(\myminixbar/_0307_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0386_ ) );
NOR2_X1 \myminixbar/_0791_ ( .A1(\myminixbar/_0309_ ), .A2(\myminixbar/_0323_ ), .ZN(\myminixbar/_0387_ ) );
BUF_X4 \myminixbar/_0792_ ( .A(\myminixbar/_0201_ ), .Z(\myminixbar/_0324_ ) );
NOR2_X1 \myminixbar/_0793_ ( .A1(\myminixbar/_0311_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0388_ ) );
NOR2_X1 \myminixbar/_0794_ ( .A1(\myminixbar/_0315_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0389_ ) );
NOR2_X1 \myminixbar/_0795_ ( .A1(\myminixbar/_0317_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0390_ ) );
NOR2_X1 \myminixbar/_0796_ ( .A1(\myminixbar/_0319_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0392_ ) );
NOR2_X1 \myminixbar/_0797_ ( .A1(\myminixbar/_0321_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0393_ ) );
AND2_X1 \myminixbar/_0798_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0495_ ), .ZN(\myminixbar/_0325_ ) );
AOI21_X2 \myminixbar/_0799_ ( .A(\myminixbar/_0325_ ), .B1(\myminixbar/_0497_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0326_ ) );
NOR2_X1 \myminixbar/_0800_ ( .A1(\myminixbar/_0326_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0491_ ) );
AND2_X1 \myminixbar/_0801_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0496_ ), .ZN(\myminixbar/_0327_ ) );
AOI21_X2 \myminixbar/_0802_ ( .A(\myminixbar/_0327_ ), .B1(\myminixbar/_0498_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0328_ ) );
NOR2_X1 \myminixbar/_0803_ ( .A1(\myminixbar/_0328_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0492_ ) );
NOR2_X1 \myminixbar/_0804_ ( .A1(\myminixbar/_0326_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0493_ ) );
NOR2_X1 \myminixbar/_0805_ ( .A1(\myminixbar/_0328_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0494_ ) );
NOR2_X1 \myminixbar/_0806_ ( .A1(\myminixbar/_0197_ ), .A2(\myminixbar/_0209_ ), .ZN(\myminixbar/_0490_ ) );
AND2_X1 \myminixbar/_0807_ ( .A1(\myminixbar/_0305_ ), .A2(\myminixbar/_0473_ ), .ZN(\myminixbar/_0329_ ) );
AOI21_X2 \myminixbar/_0808_ ( .A(\myminixbar/_0329_ ), .B1(\myminixbar/_0477_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0330_ ) );
NOR2_X1 \myminixbar/_0809_ ( .A1(\myminixbar/_0330_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0465_ ) );
AND2_X1 \myminixbar/_0810_ ( .A1(\myminixbar/_0196_ ), .A2(\myminixbar/_0474_ ), .ZN(\myminixbar/_0331_ ) );
AOI21_X1 \myminixbar/_0811_ ( .A(\myminixbar/_0331_ ), .B1(\myminixbar/_0478_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0332_ ) );
NOR2_X1 \myminixbar/_0812_ ( .A1(\myminixbar/_0332_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0466_ ) );
AND2_X1 \myminixbar/_0813_ ( .A1(\myminixbar/_0196_ ), .A2(\myminixbar/_0475_ ), .ZN(\myminixbar/_0333_ ) );
AOI21_X1 \myminixbar/_0814_ ( .A(\myminixbar/_0333_ ), .B1(\myminixbar/_0479_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0334_ ) );
NOR2_X1 \myminixbar/_0815_ ( .A1(\myminixbar/_0334_ ), .A2(\myminixbar/_0312_ ), .ZN(\myminixbar/_0467_ ) );
AND2_X1 \myminixbar/_0816_ ( .A1(\myminixbar/_0196_ ), .A2(\myminixbar/_0476_ ), .ZN(\myminixbar/_0335_ ) );
AOI21_X1 \myminixbar/_0817_ ( .A(\myminixbar/_0335_ ), .B1(\myminixbar/_0480_ ), .B2(\myminixbar/_0314_ ), .ZN(\myminixbar/_0336_ ) );
NOR2_X1 \myminixbar/_0818_ ( .A1(\myminixbar/_0336_ ), .A2(\myminixbar/_0199_ ), .ZN(\myminixbar/_0468_ ) );
NOR2_X1 \myminixbar/_0819_ ( .A1(\myminixbar/_0330_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0469_ ) );
NOR2_X1 \myminixbar/_0820_ ( .A1(\myminixbar/_0332_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0470_ ) );
NOR2_X1 \myminixbar/_0821_ ( .A1(\myminixbar/_0334_ ), .A2(\myminixbar/_0324_ ), .ZN(\myminixbar/_0471_ ) );
NOR2_X1 \myminixbar/_0822_ ( .A1(\myminixbar/_0336_ ), .A2(\myminixbar/_0201_ ), .ZN(\myminixbar/_0472_ ) );
DFF_X1 \myminixbar/_0823_ ( .D(\myminixbar/_0000_ ), .CK(clock ), .Q(\myminixbar/state [0] ), .QN(\myminixbar/_0507_ ) );
DFF_X1 \myminixbar/_0824_ ( .D(\myminixbar/_0001_ ), .CK(clock ), .Q(\myminixbar/state [2] ), .QN(\myminixbar/_0506_ ) );
BUF_X1 \myminixbar/_0825_ ( .A(\araddr_clint [0] ), .Z(\io_master_araddr [0] ) );
BUF_X1 \myminixbar/_0826_ ( .A(\araddr_clint [1] ), .Z(\io_master_araddr [1] ) );
BUF_X1 \myminixbar/_0827_ ( .A(\araddr_clint [2] ), .Z(\io_master_araddr [2] ) );
BUF_X1 \myminixbar/_0828_ ( .A(\araddr_clint [3] ), .Z(\io_master_araddr [3] ) );
BUF_X1 \myminixbar/_0829_ ( .A(\araddr_clint [4] ), .Z(\io_master_araddr [4] ) );
BUF_X1 \myminixbar/_0830_ ( .A(\araddr_clint [5] ), .Z(\io_master_araddr [5] ) );
BUF_X1 \myminixbar/_0831_ ( .A(\araddr_clint [6] ), .Z(\io_master_araddr [6] ) );
BUF_X1 \myminixbar/_0832_ ( .A(\araddr_clint [7] ), .Z(\io_master_araddr [7] ) );
BUF_X1 \myminixbar/_0833_ ( .A(\araddr_clint [8] ), .Z(\io_master_araddr [8] ) );
BUF_X1 \myminixbar/_0834_ ( .A(\araddr_clint [9] ), .Z(\io_master_araddr [9] ) );
BUF_X1 \myminixbar/_0835_ ( .A(\araddr_clint [10] ), .Z(\io_master_araddr [10] ) );
BUF_X1 \myminixbar/_0836_ ( .A(\araddr_clint [11] ), .Z(\io_master_araddr [11] ) );
BUF_X1 \myminixbar/_0837_ ( .A(\araddr_clint [12] ), .Z(\io_master_araddr [12] ) );
BUF_X1 \myminixbar/_0838_ ( .A(\araddr_clint [13] ), .Z(\io_master_araddr [13] ) );
BUF_X1 \myminixbar/_0839_ ( .A(\araddr_clint [14] ), .Z(\io_master_araddr [14] ) );
BUF_X1 \myminixbar/_0840_ ( .A(\araddr_clint [15] ), .Z(\io_master_araddr [15] ) );
BUF_X1 \myminixbar/_0841_ ( .A(\araddr_clint [16] ), .Z(\io_master_araddr [16] ) );
BUF_X1 \myminixbar/_0842_ ( .A(\araddr_clint [17] ), .Z(\io_master_araddr [17] ) );
BUF_X1 \myminixbar/_0843_ ( .A(\araddr_clint [18] ), .Z(\io_master_araddr [18] ) );
BUF_X1 \myminixbar/_0844_ ( .A(\araddr_clint [19] ), .Z(\io_master_araddr [19] ) );
BUF_X1 \myminixbar/_0845_ ( .A(\araddr_clint [20] ), .Z(\io_master_araddr [20] ) );
BUF_X1 \myminixbar/_0846_ ( .A(\araddr_clint [21] ), .Z(\io_master_araddr [21] ) );
BUF_X1 \myminixbar/_0847_ ( .A(\araddr_clint [22] ), .Z(\io_master_araddr [22] ) );
BUF_X1 \myminixbar/_0848_ ( .A(\araddr_clint [23] ), .Z(\io_master_araddr [23] ) );
BUF_X1 \myminixbar/_0849_ ( .A(\araddr_clint [24] ), .Z(\io_master_araddr [24] ) );
BUF_X1 \myminixbar/_0850_ ( .A(\araddr_clint [25] ), .Z(\io_master_araddr [25] ) );
BUF_X1 \myminixbar/_0851_ ( .A(\araddr_clint [26] ), .Z(\io_master_araddr [26] ) );
BUF_X1 \myminixbar/_0852_ ( .A(\araddr_clint [27] ), .Z(\io_master_araddr [27] ) );
BUF_X1 \myminixbar/_0853_ ( .A(\araddr_clint [28] ), .Z(\io_master_araddr [28] ) );
BUF_X1 \myminixbar/_0854_ ( .A(\araddr_clint [29] ), .Z(\io_master_araddr [29] ) );
BUF_X1 \myminixbar/_0855_ ( .A(\araddr_clint [30] ), .Z(\io_master_araddr [30] ) );
BUF_X1 \myminixbar/_0856_ ( .A(\araddr_clint [31] ), .Z(\io_master_araddr [31] ) );
BUF_X1 \myminixbar/_0857_ ( .A(\arid_clint [0] ), .Z(\io_master_arid [0] ) );
BUF_X1 \myminixbar/_0858_ ( .A(\arid_clint [1] ), .Z(\io_master_arid [1] ) );
BUF_X1 \myminixbar/_0859_ ( .A(\arid_clint [2] ), .Z(\io_master_arid [2] ) );
BUF_X1 \myminixbar/_0860_ ( .A(\arid_clint [3] ), .Z(\io_master_arid [3] ) );
BUF_X1 \myminixbar/_0861_ ( .A(\awaddr_LSU [0] ), .Z(\io_master_awaddr [0] ) );
BUF_X1 \myminixbar/_0862_ ( .A(\awaddr_LSU [1] ), .Z(\io_master_awaddr [1] ) );
BUF_X1 \myminixbar/_0863_ ( .A(\awaddr_LSU [2] ), .Z(\io_master_awaddr [2] ) );
BUF_X1 \myminixbar/_0864_ ( .A(\awaddr_LSU [3] ), .Z(\io_master_awaddr [3] ) );
BUF_X1 \myminixbar/_0865_ ( .A(\awaddr_LSU [4] ), .Z(\io_master_awaddr [4] ) );
BUF_X1 \myminixbar/_0866_ ( .A(\awaddr_LSU [5] ), .Z(\io_master_awaddr [5] ) );
BUF_X1 \myminixbar/_0867_ ( .A(\awaddr_LSU [6] ), .Z(\io_master_awaddr [6] ) );
BUF_X1 \myminixbar/_0868_ ( .A(\awaddr_LSU [7] ), .Z(\io_master_awaddr [7] ) );
BUF_X1 \myminixbar/_0869_ ( .A(\awaddr_LSU [8] ), .Z(\io_master_awaddr [8] ) );
BUF_X1 \myminixbar/_0870_ ( .A(\awaddr_LSU [9] ), .Z(\io_master_awaddr [9] ) );
BUF_X1 \myminixbar/_0871_ ( .A(\awaddr_LSU [10] ), .Z(\io_master_awaddr [10] ) );
BUF_X1 \myminixbar/_0872_ ( .A(\awaddr_LSU [11] ), .Z(\io_master_awaddr [11] ) );
BUF_X1 \myminixbar/_0873_ ( .A(\awaddr_LSU [12] ), .Z(\io_master_awaddr [12] ) );
BUF_X1 \myminixbar/_0874_ ( .A(\awaddr_LSU [13] ), .Z(\io_master_awaddr [13] ) );
BUF_X1 \myminixbar/_0875_ ( .A(\awaddr_LSU [14] ), .Z(\io_master_awaddr [14] ) );
BUF_X1 \myminixbar/_0876_ ( .A(\awaddr_LSU [15] ), .Z(\io_master_awaddr [15] ) );
BUF_X1 \myminixbar/_0877_ ( .A(\awaddr_LSU [16] ), .Z(\io_master_awaddr [16] ) );
BUF_X1 \myminixbar/_0878_ ( .A(\awaddr_LSU [17] ), .Z(\io_master_awaddr [17] ) );
BUF_X1 \myminixbar/_0879_ ( .A(\awaddr_LSU [18] ), .Z(\io_master_awaddr [18] ) );
BUF_X1 \myminixbar/_0880_ ( .A(\awaddr_LSU [19] ), .Z(\io_master_awaddr [19] ) );
BUF_X1 \myminixbar/_0881_ ( .A(\awaddr_LSU [20] ), .Z(\io_master_awaddr [20] ) );
BUF_X1 \myminixbar/_0882_ ( .A(\awaddr_LSU [21] ), .Z(\io_master_awaddr [21] ) );
BUF_X1 \myminixbar/_0883_ ( .A(\awaddr_LSU [22] ), .Z(\io_master_awaddr [22] ) );
BUF_X1 \myminixbar/_0884_ ( .A(\awaddr_LSU [23] ), .Z(\io_master_awaddr [23] ) );
BUF_X1 \myminixbar/_0885_ ( .A(\awaddr_LSU [24] ), .Z(\io_master_awaddr [24] ) );
BUF_X1 \myminixbar/_0886_ ( .A(\awaddr_LSU [25] ), .Z(\io_master_awaddr [25] ) );
BUF_X1 \myminixbar/_0887_ ( .A(\awaddr_LSU [26] ), .Z(\io_master_awaddr [26] ) );
BUF_X1 \myminixbar/_0888_ ( .A(\awaddr_LSU [27] ), .Z(\io_master_awaddr [27] ) );
BUF_X1 \myminixbar/_0889_ ( .A(\awaddr_LSU [28] ), .Z(\io_master_awaddr [28] ) );
BUF_X1 \myminixbar/_0890_ ( .A(\awaddr_LSU [29] ), .Z(\io_master_awaddr [29] ) );
BUF_X1 \myminixbar/_0891_ ( .A(\awaddr_LSU [30] ), .Z(\io_master_awaddr [30] ) );
BUF_X1 \myminixbar/_0892_ ( .A(\awaddr_LSU [31] ), .Z(\io_master_awaddr [31] ) );
BUF_X1 \myminixbar/_0893_ ( .A(\awburst_LSU [0] ), .Z(\io_master_awburst [0] ) );
BUF_X1 \myminixbar/_0894_ ( .A(\awburst_LSU [1] ), .Z(\io_master_awburst [1] ) );
BUF_X1 \myminixbar/_0895_ ( .A(\awid_LSU [0] ), .Z(\io_master_awid [0] ) );
BUF_X1 \myminixbar/_0896_ ( .A(\awid_LSU [1] ), .Z(\io_master_awid [1] ) );
BUF_X1 \myminixbar/_0897_ ( .A(\awid_LSU [2] ), .Z(\io_master_awid [2] ) );
BUF_X1 \myminixbar/_0898_ ( .A(\awid_LSU [3] ), .Z(\io_master_awid [3] ) );
BUF_X1 \myminixbar/_0899_ ( .A(\awlen_LSU [0] ), .Z(\io_master_awlen [0] ) );
BUF_X1 \myminixbar/_0900_ ( .A(\awlen_LSU [1] ), .Z(\io_master_awlen [1] ) );
BUF_X1 \myminixbar/_0901_ ( .A(\awlen_LSU [2] ), .Z(\io_master_awlen [2] ) );
BUF_X1 \myminixbar/_0902_ ( .A(\awlen_LSU [3] ), .Z(\io_master_awlen [3] ) );
BUF_X1 \myminixbar/_0903_ ( .A(\awlen_LSU [4] ), .Z(\io_master_awlen [4] ) );
BUF_X1 \myminixbar/_0904_ ( .A(\awlen_LSU [5] ), .Z(\io_master_awlen [5] ) );
BUF_X1 \myminixbar/_0905_ ( .A(\awlen_LSU [6] ), .Z(\io_master_awlen [6] ) );
BUF_X1 \myminixbar/_0906_ ( .A(\awlen_LSU [7] ), .Z(\io_master_awlen [7] ) );
BUF_X1 \myminixbar/_0907_ ( .A(io_master_awready ), .Z(awready_LSU ) );
BUF_X1 \myminixbar/_0908_ ( .A(\awsize_LSU [0] ), .Z(\io_master_awsize [0] ) );
BUF_X1 \myminixbar/_0909_ ( .A(\awsize_LSU [1] ), .Z(\io_master_awsize [1] ) );
BUF_X1 \myminixbar/_0910_ ( .A(\awsize_LSU [2] ), .Z(\io_master_awsize [2] ) );
BUF_X1 \myminixbar/_0911_ ( .A(awvalid_LSU ), .Z(io_master_awvalid ) );
BUF_X1 \myminixbar/_0912_ ( .A(\io_master_bid [0] ), .Z(\bid_LSU [0] ) );
BUF_X1 \myminixbar/_0913_ ( .A(\io_master_bid [1] ), .Z(\bid_LSU [1] ) );
BUF_X1 \myminixbar/_0914_ ( .A(\io_master_bid [2] ), .Z(\bid_LSU [2] ) );
BUF_X1 \myminixbar/_0915_ ( .A(\io_master_bid [3] ), .Z(\bid_LSU [3] ) );
BUF_X1 \myminixbar/_0916_ ( .A(bready_LSU ), .Z(io_master_bready ) );
BUF_X1 \myminixbar/_0917_ ( .A(\io_master_bresp [0] ), .Z(\bresp_LSU [0] ) );
BUF_X1 \myminixbar/_0918_ ( .A(\io_master_bresp [1] ), .Z(\bresp_LSU [1] ) );
BUF_X1 \myminixbar/_0919_ ( .A(io_master_bvalid ), .Z(bvalid_LSU ) );
BUF_X1 \myminixbar/_0920_ ( .A(\wdata_LSU [0] ), .Z(\io_master_wdata [0] ) );
BUF_X1 \myminixbar/_0921_ ( .A(\wdata_LSU [1] ), .Z(\io_master_wdata [1] ) );
BUF_X1 \myminixbar/_0922_ ( .A(\wdata_LSU [2] ), .Z(\io_master_wdata [2] ) );
BUF_X1 \myminixbar/_0923_ ( .A(\wdata_LSU [3] ), .Z(\io_master_wdata [3] ) );
BUF_X1 \myminixbar/_0924_ ( .A(\wdata_LSU [4] ), .Z(\io_master_wdata [4] ) );
BUF_X1 \myminixbar/_0925_ ( .A(\wdata_LSU [5] ), .Z(\io_master_wdata [5] ) );
BUF_X1 \myminixbar/_0926_ ( .A(\wdata_LSU [6] ), .Z(\io_master_wdata [6] ) );
BUF_X1 \myminixbar/_0927_ ( .A(\wdata_LSU [7] ), .Z(\io_master_wdata [7] ) );
BUF_X1 \myminixbar/_0928_ ( .A(\wdata_LSU [8] ), .Z(\io_master_wdata [8] ) );
BUF_X1 \myminixbar/_0929_ ( .A(\wdata_LSU [9] ), .Z(\io_master_wdata [9] ) );
BUF_X1 \myminixbar/_0930_ ( .A(\wdata_LSU [10] ), .Z(\io_master_wdata [10] ) );
BUF_X1 \myminixbar/_0931_ ( .A(\wdata_LSU [11] ), .Z(\io_master_wdata [11] ) );
BUF_X1 \myminixbar/_0932_ ( .A(\wdata_LSU [12] ), .Z(\io_master_wdata [12] ) );
BUF_X1 \myminixbar/_0933_ ( .A(\wdata_LSU [13] ), .Z(\io_master_wdata [13] ) );
BUF_X1 \myminixbar/_0934_ ( .A(\wdata_LSU [14] ), .Z(\io_master_wdata [14] ) );
BUF_X1 \myminixbar/_0935_ ( .A(\wdata_LSU [15] ), .Z(\io_master_wdata [15] ) );
BUF_X1 \myminixbar/_0936_ ( .A(\wdata_LSU [16] ), .Z(\io_master_wdata [16] ) );
BUF_X1 \myminixbar/_0937_ ( .A(\wdata_LSU [17] ), .Z(\io_master_wdata [17] ) );
BUF_X1 \myminixbar/_0938_ ( .A(\wdata_LSU [18] ), .Z(\io_master_wdata [18] ) );
BUF_X1 \myminixbar/_0939_ ( .A(\wdata_LSU [19] ), .Z(\io_master_wdata [19] ) );
BUF_X1 \myminixbar/_0940_ ( .A(\wdata_LSU [20] ), .Z(\io_master_wdata [20] ) );
BUF_X1 \myminixbar/_0941_ ( .A(\wdata_LSU [21] ), .Z(\io_master_wdata [21] ) );
BUF_X1 \myminixbar/_0942_ ( .A(\wdata_LSU [22] ), .Z(\io_master_wdata [22] ) );
BUF_X1 \myminixbar/_0943_ ( .A(\wdata_LSU [23] ), .Z(\io_master_wdata [23] ) );
BUF_X1 \myminixbar/_0944_ ( .A(\wdata_LSU [24] ), .Z(\io_master_wdata [24] ) );
BUF_X1 \myminixbar/_0945_ ( .A(\wdata_LSU [25] ), .Z(\io_master_wdata [25] ) );
BUF_X1 \myminixbar/_0946_ ( .A(\wdata_LSU [26] ), .Z(\io_master_wdata [26] ) );
BUF_X1 \myminixbar/_0947_ ( .A(\wdata_LSU [27] ), .Z(\io_master_wdata [27] ) );
BUF_X1 \myminixbar/_0948_ ( .A(\wdata_LSU [28] ), .Z(\io_master_wdata [28] ) );
BUF_X1 \myminixbar/_0949_ ( .A(\wdata_LSU [29] ), .Z(\io_master_wdata [29] ) );
BUF_X1 \myminixbar/_0950_ ( .A(\wdata_LSU [30] ), .Z(\io_master_wdata [30] ) );
BUF_X1 \myminixbar/_0951_ ( .A(\wdata_LSU [31] ), .Z(\io_master_wdata [31] ) );
BUF_X1 \myminixbar/_0952_ ( .A(wlast_LSU ), .Z(io_master_wlast ) );
BUF_X1 \myminixbar/_0953_ ( .A(io_master_wready ), .Z(wready_LSU ) );
BUF_X1 \myminixbar/_0954_ ( .A(\wstrb_LSU [0] ), .Z(\io_master_wstrb [0] ) );
BUF_X1 \myminixbar/_0955_ ( .A(\wstrb_LSU [1] ), .Z(\io_master_wstrb [1] ) );
BUF_X1 \myminixbar/_0956_ ( .A(\wstrb_LSU [2] ), .Z(\io_master_wstrb [2] ) );
BUF_X1 \myminixbar/_0957_ ( .A(\wstrb_LSU [3] ), .Z(\io_master_wstrb [3] ) );
BUF_X1 \myminixbar/_0958_ ( .A(wvalid_LSU ), .Z(io_master_wvalid ) );
BUF_X1 \myminixbar/_0959_ ( .A(\araddr_IFU [25] ), .Z(\myminixbar/_0021_ ) );
BUF_X1 \myminixbar/_0960_ ( .A(\araddr_LSU [25] ), .Z(\myminixbar/_0053_ ) );
BUF_X1 \myminixbar/_0961_ ( .A(rmem_quest_LSU ), .Z(\myminixbar/_0486_ ) );
BUF_X1 \myminixbar/_0962_ ( .A(\myminixbar/state [2] ), .Z(\myminixbar/_0505_ ) );
BUF_X1 \myminixbar/_0963_ ( .A(\myminixbar/state [0] ), .Z(\myminixbar/_0504_ ) );
BUF_X1 \myminixbar/_0964_ ( .A(rmem_quest_IFU ), .Z(\myminixbar/_0485_ ) );
BUF_X1 \myminixbar/_0965_ ( .A(\myminixbar/_0085_ ), .Z(\araddr_clint [25] ) );
BUF_X1 \myminixbar/_0966_ ( .A(\araddr_LSU [16] ), .Z(\myminixbar/_0043_ ) );
BUF_X1 \myminixbar/_0967_ ( .A(\araddr_IFU [16] ), .Z(\myminixbar/_0011_ ) );
BUF_X1 \myminixbar/_0968_ ( .A(\myminixbar/_0075_ ), .Z(\araddr_clint [16] ) );
BUF_X1 \myminixbar/_0969_ ( .A(\araddr_LSU [17] ), .Z(\myminixbar/_0044_ ) );
BUF_X1 \myminixbar/_0970_ ( .A(\araddr_IFU [17] ), .Z(\myminixbar/_0012_ ) );
BUF_X1 \myminixbar/_0971_ ( .A(\myminixbar/_0076_ ), .Z(\araddr_clint [17] ) );
BUF_X1 \myminixbar/_0972_ ( .A(\araddr_LSU [18] ), .Z(\myminixbar/_0045_ ) );
BUF_X1 \myminixbar/_0973_ ( .A(\araddr_IFU [18] ), .Z(\myminixbar/_0013_ ) );
BUF_X1 \myminixbar/_0974_ ( .A(\myminixbar/_0077_ ), .Z(\araddr_clint [18] ) );
BUF_X1 \myminixbar/_0975_ ( .A(\araddr_LSU [19] ), .Z(\myminixbar/_0046_ ) );
BUF_X1 \myminixbar/_0976_ ( .A(\araddr_IFU [19] ), .Z(\myminixbar/_0014_ ) );
BUF_X1 \myminixbar/_0977_ ( .A(\myminixbar/_0078_ ), .Z(\araddr_clint [19] ) );
BUF_X1 \myminixbar/_0978_ ( .A(\araddr_LSU [20] ), .Z(\myminixbar/_0048_ ) );
BUF_X1 \myminixbar/_0979_ ( .A(\araddr_IFU [20] ), .Z(\myminixbar/_0016_ ) );
BUF_X1 \myminixbar/_0980_ ( .A(\myminixbar/_0080_ ), .Z(\araddr_clint [20] ) );
BUF_X1 \myminixbar/_0981_ ( .A(\araddr_LSU [21] ), .Z(\myminixbar/_0049_ ) );
BUF_X1 \myminixbar/_0982_ ( .A(\araddr_IFU [21] ), .Z(\myminixbar/_0017_ ) );
BUF_X1 \myminixbar/_0983_ ( .A(\myminixbar/_0081_ ), .Z(\araddr_clint [21] ) );
BUF_X1 \myminixbar/_0984_ ( .A(\araddr_LSU [22] ), .Z(\myminixbar/_0050_ ) );
BUF_X1 \myminixbar/_0985_ ( .A(\araddr_IFU [22] ), .Z(\myminixbar/_0018_ ) );
BUF_X1 \myminixbar/_0986_ ( .A(\myminixbar/_0082_ ), .Z(\araddr_clint [22] ) );
BUF_X1 \myminixbar/_0987_ ( .A(\araddr_LSU [23] ), .Z(\myminixbar/_0051_ ) );
BUF_X1 \myminixbar/_0988_ ( .A(\araddr_IFU [23] ), .Z(\myminixbar/_0019_ ) );
BUF_X1 \myminixbar/_0989_ ( .A(\myminixbar/_0083_ ), .Z(\araddr_clint [23] ) );
BUF_X1 \myminixbar/_0990_ ( .A(\araddr_LSU [24] ), .Z(\myminixbar/_0052_ ) );
BUF_X1 \myminixbar/_0991_ ( .A(\araddr_IFU [24] ), .Z(\myminixbar/_0020_ ) );
BUF_X1 \myminixbar/_0992_ ( .A(\myminixbar/_0084_ ), .Z(\araddr_clint [24] ) );
BUF_X1 \myminixbar/_0993_ ( .A(\araddr_LSU [26] ), .Z(\myminixbar/_0054_ ) );
BUF_X1 \myminixbar/_0994_ ( .A(\araddr_IFU [26] ), .Z(\myminixbar/_0022_ ) );
BUF_X1 \myminixbar/_0995_ ( .A(\myminixbar/_0086_ ), .Z(\araddr_clint [26] ) );
BUF_X1 \myminixbar/_0996_ ( .A(\araddr_LSU [27] ), .Z(\myminixbar/_0055_ ) );
BUF_X1 \myminixbar/_0997_ ( .A(\araddr_IFU [27] ), .Z(\myminixbar/_0023_ ) );
BUF_X1 \myminixbar/_0998_ ( .A(\myminixbar/_0087_ ), .Z(\araddr_clint [27] ) );
BUF_X1 \myminixbar/_0999_ ( .A(\araddr_LSU [28] ), .Z(\myminixbar/_0056_ ) );
BUF_X1 \myminixbar/_1000_ ( .A(\araddr_IFU [28] ), .Z(\myminixbar/_0024_ ) );
BUF_X1 \myminixbar/_1001_ ( .A(\myminixbar/_0088_ ), .Z(\araddr_clint [28] ) );
BUF_X1 \myminixbar/_1002_ ( .A(\araddr_LSU [29] ), .Z(\myminixbar/_0057_ ) );
BUF_X1 \myminixbar/_1003_ ( .A(\araddr_IFU [29] ), .Z(\myminixbar/_0025_ ) );
BUF_X1 \myminixbar/_1004_ ( .A(\myminixbar/_0089_ ), .Z(\araddr_clint [29] ) );
BUF_X1 \myminixbar/_1005_ ( .A(\araddr_LSU [30] ), .Z(\myminixbar/_0059_ ) );
BUF_X1 \myminixbar/_1006_ ( .A(\araddr_IFU [30] ), .Z(\myminixbar/_0027_ ) );
BUF_X1 \myminixbar/_1007_ ( .A(\myminixbar/_0091_ ), .Z(\araddr_clint [30] ) );
BUF_X1 \myminixbar/_1008_ ( .A(\araddr_LSU [31] ), .Z(\myminixbar/_0060_ ) );
BUF_X1 \myminixbar/_1009_ ( .A(\araddr_IFU [31] ), .Z(\myminixbar/_0028_ ) );
BUF_X1 \myminixbar/_1010_ ( .A(\myminixbar/_0092_ ), .Z(\araddr_clint [31] ) );
BUF_X1 \myminixbar/_1011_ ( .A(arvalid_IFU ), .Z(\myminixbar/_0155_ ) );
BUF_X1 \myminixbar/_1012_ ( .A(arvalid_LSU ), .Z(\myminixbar/_0156_ ) );
BUF_X1 \myminixbar/_1013_ ( .A(\myminixbar/_0157_ ), .Z(arvalid_clint ) );
BUF_X1 \myminixbar/_1014_ ( .A(io_master_arready ), .Z(\myminixbar/_0145_ ) );
BUF_X1 \myminixbar/_1015_ ( .A(arready_clint ), .Z(\myminixbar/_0144_ ) );
BUF_X1 \myminixbar/_1016_ ( .A(\myminixbar/_0142_ ), .Z(arready_IFU ) );
BUF_X1 \myminixbar/_1017_ ( .A(\myminixbar/_0143_ ), .Z(arready_LSU ) );
BUF_X1 \myminixbar/_1018_ ( .A(rvalid_clint ), .Z(\myminixbar/_0502_ ) );
BUF_X1 \myminixbar/_1019_ ( .A(io_master_rvalid ), .Z(\myminixbar/_0503_ ) );
BUF_X1 \myminixbar/_1020_ ( .A(\myminixbar/_0500_ ), .Z(rvalid_IFU ) );
BUF_X1 \myminixbar/_1021_ ( .A(\myminixbar/_0501_ ), .Z(rvalid_LSU ) );
BUF_X1 \myminixbar/_1022_ ( .A(rready_IFU ), .Z(\myminixbar/_0487_ ) );
BUF_X1 \myminixbar/_1023_ ( .A(rready_LSU ), .Z(\myminixbar/_0488_ ) );
BUF_X1 \myminixbar/_1024_ ( .A(\myminixbar/_0489_ ), .Z(rready_clint ) );
BUF_X1 \myminixbar/_1025_ ( .A(rlast_clint ), .Z(\myminixbar/_0483_ ) );
BUF_X1 \myminixbar/_1026_ ( .A(io_master_rlast ), .Z(\myminixbar/_0484_ ) );
BUF_X1 \myminixbar/_1027_ ( .A(\myminixbar/_0481_ ), .Z(rlast_IFU ) );
BUF_X1 \myminixbar/_1028_ ( .A(\myminixbar/_0482_ ), .Z(rlast_LSU ) );
BUF_X1 \myminixbar/_1029_ ( .A(reset ), .Z(\myminixbar/_0499_ ) );
BUF_X1 \myminixbar/_1030_ ( .A(\myminixbar/_0002_ ), .Z(\myminixbar/_0000_ ) );
BUF_X1 \myminixbar/_1031_ ( .A(\myminixbar/_0003_ ), .Z(\myminixbar/_0001_ ) );
BUF_X1 \myminixbar/_1032_ ( .A(\araddr_LSU [0] ), .Z(\myminixbar/_0036_ ) );
BUF_X1 \myminixbar/_1033_ ( .A(\araddr_IFU [0] ), .Z(\myminixbar/_0004_ ) );
BUF_X1 \myminixbar/_1034_ ( .A(\myminixbar/_0068_ ), .Z(\araddr_clint [0] ) );
BUF_X1 \myminixbar/_1035_ ( .A(\araddr_LSU [1] ), .Z(\myminixbar/_0047_ ) );
BUF_X1 \myminixbar/_1036_ ( .A(\araddr_IFU [1] ), .Z(\myminixbar/_0015_ ) );
BUF_X1 \myminixbar/_1037_ ( .A(\myminixbar/_0079_ ), .Z(\araddr_clint [1] ) );
BUF_X1 \myminixbar/_1038_ ( .A(\araddr_LSU [2] ), .Z(\myminixbar/_0058_ ) );
BUF_X1 \myminixbar/_1039_ ( .A(\araddr_IFU [2] ), .Z(\myminixbar/_0026_ ) );
BUF_X1 \myminixbar/_1040_ ( .A(\myminixbar/_0090_ ), .Z(\araddr_clint [2] ) );
BUF_X1 \myminixbar/_1041_ ( .A(\araddr_LSU [3] ), .Z(\myminixbar/_0061_ ) );
BUF_X1 \myminixbar/_1042_ ( .A(\araddr_IFU [3] ), .Z(\myminixbar/_0029_ ) );
BUF_X1 \myminixbar/_1043_ ( .A(\myminixbar/_0093_ ), .Z(\araddr_clint [3] ) );
BUF_X1 \myminixbar/_1044_ ( .A(\araddr_LSU [4] ), .Z(\myminixbar/_0062_ ) );
BUF_X1 \myminixbar/_1045_ ( .A(\araddr_IFU [4] ), .Z(\myminixbar/_0030_ ) );
BUF_X1 \myminixbar/_1046_ ( .A(\myminixbar/_0094_ ), .Z(\araddr_clint [4] ) );
BUF_X1 \myminixbar/_1047_ ( .A(\araddr_LSU [5] ), .Z(\myminixbar/_0063_ ) );
BUF_X1 \myminixbar/_1048_ ( .A(\araddr_IFU [5] ), .Z(\myminixbar/_0031_ ) );
BUF_X1 \myminixbar/_1049_ ( .A(\myminixbar/_0095_ ), .Z(\araddr_clint [5] ) );
BUF_X1 \myminixbar/_1050_ ( .A(\araddr_LSU [6] ), .Z(\myminixbar/_0064_ ) );
BUF_X1 \myminixbar/_1051_ ( .A(\araddr_IFU [6] ), .Z(\myminixbar/_0032_ ) );
BUF_X1 \myminixbar/_1052_ ( .A(\myminixbar/_0096_ ), .Z(\araddr_clint [6] ) );
BUF_X1 \myminixbar/_1053_ ( .A(\araddr_LSU [7] ), .Z(\myminixbar/_0065_ ) );
BUF_X1 \myminixbar/_1054_ ( .A(\araddr_IFU [7] ), .Z(\myminixbar/_0033_ ) );
BUF_X1 \myminixbar/_1055_ ( .A(\myminixbar/_0097_ ), .Z(\araddr_clint [7] ) );
BUF_X1 \myminixbar/_1056_ ( .A(\araddr_LSU [8] ), .Z(\myminixbar/_0066_ ) );
BUF_X1 \myminixbar/_1057_ ( .A(\araddr_IFU [8] ), .Z(\myminixbar/_0034_ ) );
BUF_X1 \myminixbar/_1058_ ( .A(\myminixbar/_0098_ ), .Z(\araddr_clint [8] ) );
BUF_X1 \myminixbar/_1059_ ( .A(\araddr_LSU [9] ), .Z(\myminixbar/_0067_ ) );
BUF_X1 \myminixbar/_1060_ ( .A(\araddr_IFU [9] ), .Z(\myminixbar/_0035_ ) );
BUF_X1 \myminixbar/_1061_ ( .A(\myminixbar/_0099_ ), .Z(\araddr_clint [9] ) );
BUF_X1 \myminixbar/_1062_ ( .A(\araddr_LSU [10] ), .Z(\myminixbar/_0037_ ) );
BUF_X1 \myminixbar/_1063_ ( .A(\araddr_IFU [10] ), .Z(\myminixbar/_0005_ ) );
BUF_X1 \myminixbar/_1064_ ( .A(\myminixbar/_0069_ ), .Z(\araddr_clint [10] ) );
BUF_X1 \myminixbar/_1065_ ( .A(\araddr_LSU [11] ), .Z(\myminixbar/_0038_ ) );
BUF_X1 \myminixbar/_1066_ ( .A(\araddr_IFU [11] ), .Z(\myminixbar/_0006_ ) );
BUF_X1 \myminixbar/_1067_ ( .A(\myminixbar/_0070_ ), .Z(\araddr_clint [11] ) );
BUF_X1 \myminixbar/_1068_ ( .A(\araddr_LSU [12] ), .Z(\myminixbar/_0039_ ) );
BUF_X1 \myminixbar/_1069_ ( .A(\araddr_IFU [12] ), .Z(\myminixbar/_0007_ ) );
BUF_X1 \myminixbar/_1070_ ( .A(\myminixbar/_0071_ ), .Z(\araddr_clint [12] ) );
BUF_X1 \myminixbar/_1071_ ( .A(\araddr_LSU [13] ), .Z(\myminixbar/_0040_ ) );
BUF_X1 \myminixbar/_1072_ ( .A(\araddr_IFU [13] ), .Z(\myminixbar/_0008_ ) );
BUF_X1 \myminixbar/_1073_ ( .A(\myminixbar/_0072_ ), .Z(\araddr_clint [13] ) );
BUF_X1 \myminixbar/_1074_ ( .A(\araddr_LSU [14] ), .Z(\myminixbar/_0041_ ) );
BUF_X1 \myminixbar/_1075_ ( .A(\araddr_IFU [14] ), .Z(\myminixbar/_0009_ ) );
BUF_X1 \myminixbar/_1076_ ( .A(\myminixbar/_0073_ ), .Z(\araddr_clint [14] ) );
BUF_X1 \myminixbar/_1077_ ( .A(\araddr_LSU [15] ), .Z(\myminixbar/_0042_ ) );
BUF_X1 \myminixbar/_1078_ ( .A(\araddr_IFU [15] ), .Z(\myminixbar/_0010_ ) );
BUF_X1 \myminixbar/_1079_ ( .A(\myminixbar/_0074_ ), .Z(\araddr_clint [15] ) );
BUF_X1 \myminixbar/_1080_ ( .A(\myminixbar/_0158_ ), .Z(io_master_arvalid ) );
BUF_X1 \myminixbar/_1081_ ( .A(\arid_LSU [0] ), .Z(\myminixbar/_0110_ ) );
BUF_X1 \myminixbar/_1082_ ( .A(\arid_IFU [0] ), .Z(\myminixbar/_0106_ ) );
BUF_X1 \myminixbar/_1083_ ( .A(\myminixbar/_0114_ ), .Z(\arid_clint [0] ) );
BUF_X1 \myminixbar/_1084_ ( .A(\arid_LSU [1] ), .Z(\myminixbar/_0111_ ) );
BUF_X1 \myminixbar/_1085_ ( .A(\arid_IFU [1] ), .Z(\myminixbar/_0107_ ) );
BUF_X1 \myminixbar/_1086_ ( .A(\myminixbar/_0115_ ), .Z(\arid_clint [1] ) );
BUF_X1 \myminixbar/_1087_ ( .A(\arid_LSU [2] ), .Z(\myminixbar/_0112_ ) );
BUF_X1 \myminixbar/_1088_ ( .A(\arid_IFU [2] ), .Z(\myminixbar/_0108_ ) );
BUF_X1 \myminixbar/_1089_ ( .A(\myminixbar/_0116_ ), .Z(\arid_clint [2] ) );
BUF_X1 \myminixbar/_1090_ ( .A(\arid_LSU [3] ), .Z(\myminixbar/_0113_ ) );
BUF_X1 \myminixbar/_1091_ ( .A(\arid_IFU [3] ), .Z(\myminixbar/_0109_ ) );
BUF_X1 \myminixbar/_1092_ ( .A(\myminixbar/_0117_ ), .Z(\arid_clint [3] ) );
BUF_X1 \myminixbar/_1093_ ( .A(\arlen_LSU [0] ), .Z(\myminixbar/_0126_ ) );
BUF_X1 \myminixbar/_1094_ ( .A(\arlen_IFU [0] ), .Z(\myminixbar/_0118_ ) );
BUF_X1 \myminixbar/_1095_ ( .A(\myminixbar/_0134_ ), .Z(\io_master_arlen [0] ) );
BUF_X1 \myminixbar/_1096_ ( .A(\arlen_LSU [1] ), .Z(\myminixbar/_0127_ ) );
BUF_X1 \myminixbar/_1097_ ( .A(\arlen_IFU [1] ), .Z(\myminixbar/_0119_ ) );
BUF_X1 \myminixbar/_1098_ ( .A(\myminixbar/_0135_ ), .Z(\io_master_arlen [1] ) );
BUF_X1 \myminixbar/_1099_ ( .A(\arlen_LSU [2] ), .Z(\myminixbar/_0128_ ) );
BUF_X1 \myminixbar/_1100_ ( .A(\arlen_IFU [2] ), .Z(\myminixbar/_0120_ ) );
BUF_X1 \myminixbar/_1101_ ( .A(\myminixbar/_0136_ ), .Z(\io_master_arlen [2] ) );
BUF_X1 \myminixbar/_1102_ ( .A(\arlen_LSU [3] ), .Z(\myminixbar/_0129_ ) );
BUF_X1 \myminixbar/_1103_ ( .A(\arlen_IFU [3] ), .Z(\myminixbar/_0121_ ) );
BUF_X1 \myminixbar/_1104_ ( .A(\myminixbar/_0137_ ), .Z(\io_master_arlen [3] ) );
BUF_X1 \myminixbar/_1105_ ( .A(\arlen_LSU [4] ), .Z(\myminixbar/_0130_ ) );
BUF_X1 \myminixbar/_1106_ ( .A(\arlen_IFU [4] ), .Z(\myminixbar/_0122_ ) );
BUF_X1 \myminixbar/_1107_ ( .A(\myminixbar/_0138_ ), .Z(\io_master_arlen [4] ) );
BUF_X1 \myminixbar/_1108_ ( .A(\arlen_LSU [5] ), .Z(\myminixbar/_0131_ ) );
BUF_X1 \myminixbar/_1109_ ( .A(\arlen_IFU [5] ), .Z(\myminixbar/_0123_ ) );
BUF_X1 \myminixbar/_1110_ ( .A(\myminixbar/_0139_ ), .Z(\io_master_arlen [5] ) );
BUF_X1 \myminixbar/_1111_ ( .A(\arlen_LSU [6] ), .Z(\myminixbar/_0132_ ) );
BUF_X1 \myminixbar/_1112_ ( .A(\arlen_IFU [6] ), .Z(\myminixbar/_0124_ ) );
BUF_X1 \myminixbar/_1113_ ( .A(\myminixbar/_0140_ ), .Z(\io_master_arlen [6] ) );
BUF_X1 \myminixbar/_1114_ ( .A(\arlen_LSU [7] ), .Z(\myminixbar/_0133_ ) );
BUF_X1 \myminixbar/_1115_ ( .A(\arlen_IFU [7] ), .Z(\myminixbar/_0125_ ) );
BUF_X1 \myminixbar/_1116_ ( .A(\myminixbar/_0141_ ), .Z(\io_master_arlen [7] ) );
BUF_X1 \myminixbar/_1117_ ( .A(\arsize_LSU [0] ), .Z(\myminixbar/_0149_ ) );
BUF_X1 \myminixbar/_1118_ ( .A(\arsize_IFU [0] ), .Z(\myminixbar/_0146_ ) );
BUF_X1 \myminixbar/_1119_ ( .A(\myminixbar/_0152_ ), .Z(\io_master_arsize [0] ) );
BUF_X1 \myminixbar/_1120_ ( .A(\arsize_LSU [1] ), .Z(\myminixbar/_0150_ ) );
BUF_X1 \myminixbar/_1121_ ( .A(\arsize_IFU [1] ), .Z(\myminixbar/_0147_ ) );
BUF_X1 \myminixbar/_1122_ ( .A(\myminixbar/_0153_ ), .Z(\io_master_arsize [1] ) );
BUF_X1 \myminixbar/_1123_ ( .A(\arsize_LSU [2] ), .Z(\myminixbar/_0151_ ) );
BUF_X1 \myminixbar/_1124_ ( .A(\arsize_IFU [2] ), .Z(\myminixbar/_0148_ ) );
BUF_X1 \myminixbar/_1125_ ( .A(\myminixbar/_0154_ ), .Z(\io_master_arsize [2] ) );
BUF_X1 \myminixbar/_1126_ ( .A(\arburst_LSU [0] ), .Z(\myminixbar/_0102_ ) );
BUF_X1 \myminixbar/_1127_ ( .A(\arburst_IFU [0] ), .Z(\myminixbar/_0100_ ) );
BUF_X1 \myminixbar/_1128_ ( .A(\myminixbar/_0104_ ), .Z(\io_master_arburst [0] ) );
BUF_X1 \myminixbar/_1129_ ( .A(\arburst_LSU [1] ), .Z(\myminixbar/_0103_ ) );
BUF_X1 \myminixbar/_1130_ ( .A(\arburst_IFU [1] ), .Z(\myminixbar/_0101_ ) );
BUF_X1 \myminixbar/_1131_ ( .A(\myminixbar/_0105_ ), .Z(\io_master_arburst [1] ) );
BUF_X1 \myminixbar/_1132_ ( .A(\rdata_clint [0] ), .Z(\myminixbar/_0401_ ) );
BUF_X1 \myminixbar/_1133_ ( .A(\io_master_rdata [0] ), .Z(\myminixbar/_0433_ ) );
BUF_X1 \myminixbar/_1134_ ( .A(\myminixbar/_0337_ ), .Z(\rdata_IFU [0] ) );
BUF_X1 \myminixbar/_1135_ ( .A(\rdata_clint [1] ), .Z(\myminixbar/_0412_ ) );
BUF_X1 \myminixbar/_1136_ ( .A(\io_master_rdata [1] ), .Z(\myminixbar/_0444_ ) );
BUF_X1 \myminixbar/_1137_ ( .A(\myminixbar/_0348_ ), .Z(\rdata_IFU [1] ) );
BUF_X1 \myminixbar/_1138_ ( .A(\rdata_clint [2] ), .Z(\myminixbar/_0423_ ) );
BUF_X1 \myminixbar/_1139_ ( .A(\io_master_rdata [2] ), .Z(\myminixbar/_0455_ ) );
BUF_X1 \myminixbar/_1140_ ( .A(\myminixbar/_0359_ ), .Z(\rdata_IFU [2] ) );
BUF_X1 \myminixbar/_1141_ ( .A(\rdata_clint [3] ), .Z(\myminixbar/_0426_ ) );
BUF_X1 \myminixbar/_1142_ ( .A(\io_master_rdata [3] ), .Z(\myminixbar/_0458_ ) );
BUF_X1 \myminixbar/_1143_ ( .A(\myminixbar/_0362_ ), .Z(\rdata_IFU [3] ) );
BUF_X1 \myminixbar/_1144_ ( .A(\rdata_clint [4] ), .Z(\myminixbar/_0427_ ) );
BUF_X1 \myminixbar/_1145_ ( .A(\io_master_rdata [4] ), .Z(\myminixbar/_0459_ ) );
BUF_X1 \myminixbar/_1146_ ( .A(\myminixbar/_0363_ ), .Z(\rdata_IFU [4] ) );
BUF_X1 \myminixbar/_1147_ ( .A(\rdata_clint [5] ), .Z(\myminixbar/_0428_ ) );
BUF_X1 \myminixbar/_1148_ ( .A(\io_master_rdata [5] ), .Z(\myminixbar/_0460_ ) );
BUF_X1 \myminixbar/_1149_ ( .A(\myminixbar/_0364_ ), .Z(\rdata_IFU [5] ) );
BUF_X1 \myminixbar/_1150_ ( .A(\rdata_clint [6] ), .Z(\myminixbar/_0429_ ) );
BUF_X1 \myminixbar/_1151_ ( .A(\io_master_rdata [6] ), .Z(\myminixbar/_0461_ ) );
BUF_X1 \myminixbar/_1152_ ( .A(\myminixbar/_0365_ ), .Z(\rdata_IFU [6] ) );
BUF_X1 \myminixbar/_1153_ ( .A(\rdata_clint [7] ), .Z(\myminixbar/_0430_ ) );
BUF_X1 \myminixbar/_1154_ ( .A(\io_master_rdata [7] ), .Z(\myminixbar/_0462_ ) );
BUF_X1 \myminixbar/_1155_ ( .A(\myminixbar/_0366_ ), .Z(\rdata_IFU [7] ) );
BUF_X1 \myminixbar/_1156_ ( .A(\rdata_clint [8] ), .Z(\myminixbar/_0431_ ) );
BUF_X1 \myminixbar/_1157_ ( .A(\io_master_rdata [8] ), .Z(\myminixbar/_0463_ ) );
BUF_X1 \myminixbar/_1158_ ( .A(\myminixbar/_0367_ ), .Z(\rdata_IFU [8] ) );
BUF_X1 \myminixbar/_1159_ ( .A(\rdata_clint [9] ), .Z(\myminixbar/_0432_ ) );
BUF_X1 \myminixbar/_1160_ ( .A(\io_master_rdata [9] ), .Z(\myminixbar/_0464_ ) );
BUF_X1 \myminixbar/_1161_ ( .A(\myminixbar/_0368_ ), .Z(\rdata_IFU [9] ) );
BUF_X1 \myminixbar/_1162_ ( .A(\rdata_clint [10] ), .Z(\myminixbar/_0402_ ) );
BUF_X1 \myminixbar/_1163_ ( .A(\io_master_rdata [10] ), .Z(\myminixbar/_0434_ ) );
BUF_X1 \myminixbar/_1164_ ( .A(\myminixbar/_0338_ ), .Z(\rdata_IFU [10] ) );
BUF_X1 \myminixbar/_1165_ ( .A(\rdata_clint [11] ), .Z(\myminixbar/_0403_ ) );
BUF_X1 \myminixbar/_1166_ ( .A(\io_master_rdata [11] ), .Z(\myminixbar/_0435_ ) );
BUF_X1 \myminixbar/_1167_ ( .A(\myminixbar/_0339_ ), .Z(\rdata_IFU [11] ) );
BUF_X1 \myminixbar/_1168_ ( .A(\rdata_clint [12] ), .Z(\myminixbar/_0404_ ) );
BUF_X1 \myminixbar/_1169_ ( .A(\io_master_rdata [12] ), .Z(\myminixbar/_0436_ ) );
BUF_X1 \myminixbar/_1170_ ( .A(\myminixbar/_0340_ ), .Z(\rdata_IFU [12] ) );
BUF_X1 \myminixbar/_1171_ ( .A(\rdata_clint [13] ), .Z(\myminixbar/_0405_ ) );
BUF_X1 \myminixbar/_1172_ ( .A(\io_master_rdata [13] ), .Z(\myminixbar/_0437_ ) );
BUF_X1 \myminixbar/_1173_ ( .A(\myminixbar/_0341_ ), .Z(\rdata_IFU [13] ) );
BUF_X1 \myminixbar/_1174_ ( .A(\rdata_clint [14] ), .Z(\myminixbar/_0406_ ) );
BUF_X1 \myminixbar/_1175_ ( .A(\io_master_rdata [14] ), .Z(\myminixbar/_0438_ ) );
BUF_X1 \myminixbar/_1176_ ( .A(\myminixbar/_0342_ ), .Z(\rdata_IFU [14] ) );
BUF_X1 \myminixbar/_1177_ ( .A(\rdata_clint [15] ), .Z(\myminixbar/_0407_ ) );
BUF_X1 \myminixbar/_1178_ ( .A(\io_master_rdata [15] ), .Z(\myminixbar/_0439_ ) );
BUF_X1 \myminixbar/_1179_ ( .A(\myminixbar/_0343_ ), .Z(\rdata_IFU [15] ) );
BUF_X1 \myminixbar/_1180_ ( .A(\rdata_clint [16] ), .Z(\myminixbar/_0408_ ) );
BUF_X1 \myminixbar/_1181_ ( .A(\io_master_rdata [16] ), .Z(\myminixbar/_0440_ ) );
BUF_X1 \myminixbar/_1182_ ( .A(\myminixbar/_0344_ ), .Z(\rdata_IFU [16] ) );
BUF_X1 \myminixbar/_1183_ ( .A(\rdata_clint [17] ), .Z(\myminixbar/_0409_ ) );
BUF_X1 \myminixbar/_1184_ ( .A(\io_master_rdata [17] ), .Z(\myminixbar/_0441_ ) );
BUF_X1 \myminixbar/_1185_ ( .A(\myminixbar/_0345_ ), .Z(\rdata_IFU [17] ) );
BUF_X1 \myminixbar/_1186_ ( .A(\rdata_clint [18] ), .Z(\myminixbar/_0410_ ) );
BUF_X1 \myminixbar/_1187_ ( .A(\io_master_rdata [18] ), .Z(\myminixbar/_0442_ ) );
BUF_X1 \myminixbar/_1188_ ( .A(\myminixbar/_0346_ ), .Z(\rdata_IFU [18] ) );
BUF_X1 \myminixbar/_1189_ ( .A(\rdata_clint [19] ), .Z(\myminixbar/_0411_ ) );
BUF_X1 \myminixbar/_1190_ ( .A(\io_master_rdata [19] ), .Z(\myminixbar/_0443_ ) );
BUF_X1 \myminixbar/_1191_ ( .A(\myminixbar/_0347_ ), .Z(\rdata_IFU [19] ) );
BUF_X1 \myminixbar/_1192_ ( .A(\rdata_clint [20] ), .Z(\myminixbar/_0413_ ) );
BUF_X1 \myminixbar/_1193_ ( .A(\io_master_rdata [20] ), .Z(\myminixbar/_0445_ ) );
BUF_X1 \myminixbar/_1194_ ( .A(\myminixbar/_0349_ ), .Z(\rdata_IFU [20] ) );
BUF_X1 \myminixbar/_1195_ ( .A(\rdata_clint [21] ), .Z(\myminixbar/_0414_ ) );
BUF_X1 \myminixbar/_1196_ ( .A(\io_master_rdata [21] ), .Z(\myminixbar/_0446_ ) );
BUF_X1 \myminixbar/_1197_ ( .A(\myminixbar/_0350_ ), .Z(\rdata_IFU [21] ) );
BUF_X1 \myminixbar/_1198_ ( .A(\rdata_clint [22] ), .Z(\myminixbar/_0415_ ) );
BUF_X1 \myminixbar/_1199_ ( .A(\io_master_rdata [22] ), .Z(\myminixbar/_0447_ ) );
BUF_X1 \myminixbar/_1200_ ( .A(\myminixbar/_0351_ ), .Z(\rdata_IFU [22] ) );
BUF_X1 \myminixbar/_1201_ ( .A(\rdata_clint [23] ), .Z(\myminixbar/_0416_ ) );
BUF_X1 \myminixbar/_1202_ ( .A(\io_master_rdata [23] ), .Z(\myminixbar/_0448_ ) );
BUF_X1 \myminixbar/_1203_ ( .A(\myminixbar/_0352_ ), .Z(\rdata_IFU [23] ) );
BUF_X1 \myminixbar/_1204_ ( .A(\rdata_clint [24] ), .Z(\myminixbar/_0417_ ) );
BUF_X1 \myminixbar/_1205_ ( .A(\io_master_rdata [24] ), .Z(\myminixbar/_0449_ ) );
BUF_X1 \myminixbar/_1206_ ( .A(\myminixbar/_0353_ ), .Z(\rdata_IFU [24] ) );
BUF_X1 \myminixbar/_1207_ ( .A(\rdata_clint [25] ), .Z(\myminixbar/_0418_ ) );
BUF_X1 \myminixbar/_1208_ ( .A(\io_master_rdata [25] ), .Z(\myminixbar/_0450_ ) );
BUF_X1 \myminixbar/_1209_ ( .A(\myminixbar/_0354_ ), .Z(\rdata_IFU [25] ) );
BUF_X1 \myminixbar/_1210_ ( .A(\rdata_clint [26] ), .Z(\myminixbar/_0419_ ) );
BUF_X1 \myminixbar/_1211_ ( .A(\io_master_rdata [26] ), .Z(\myminixbar/_0451_ ) );
BUF_X1 \myminixbar/_1212_ ( .A(\myminixbar/_0355_ ), .Z(\rdata_IFU [26] ) );
BUF_X1 \myminixbar/_1213_ ( .A(\rdata_clint [27] ), .Z(\myminixbar/_0420_ ) );
BUF_X1 \myminixbar/_1214_ ( .A(\io_master_rdata [27] ), .Z(\myminixbar/_0452_ ) );
BUF_X1 \myminixbar/_1215_ ( .A(\myminixbar/_0356_ ), .Z(\rdata_IFU [27] ) );
BUF_X1 \myminixbar/_1216_ ( .A(\rdata_clint [28] ), .Z(\myminixbar/_0421_ ) );
BUF_X1 \myminixbar/_1217_ ( .A(\io_master_rdata [28] ), .Z(\myminixbar/_0453_ ) );
BUF_X1 \myminixbar/_1218_ ( .A(\myminixbar/_0357_ ), .Z(\rdata_IFU [28] ) );
BUF_X1 \myminixbar/_1219_ ( .A(\rdata_clint [29] ), .Z(\myminixbar/_0422_ ) );
BUF_X1 \myminixbar/_1220_ ( .A(\io_master_rdata [29] ), .Z(\myminixbar/_0454_ ) );
BUF_X1 \myminixbar/_1221_ ( .A(\myminixbar/_0358_ ), .Z(\rdata_IFU [29] ) );
BUF_X1 \myminixbar/_1222_ ( .A(\rdata_clint [30] ), .Z(\myminixbar/_0424_ ) );
BUF_X1 \myminixbar/_1223_ ( .A(\io_master_rdata [30] ), .Z(\myminixbar/_0456_ ) );
BUF_X1 \myminixbar/_1224_ ( .A(\myminixbar/_0360_ ), .Z(\rdata_IFU [30] ) );
BUF_X1 \myminixbar/_1225_ ( .A(\rdata_clint [31] ), .Z(\myminixbar/_0425_ ) );
BUF_X1 \myminixbar/_1226_ ( .A(\io_master_rdata [31] ), .Z(\myminixbar/_0457_ ) );
BUF_X1 \myminixbar/_1227_ ( .A(\myminixbar/_0361_ ), .Z(\rdata_IFU [31] ) );
BUF_X1 \myminixbar/_1228_ ( .A(\myminixbar/_0369_ ), .Z(\rdata_LSU [0] ) );
BUF_X1 \myminixbar/_1229_ ( .A(\myminixbar/_0380_ ), .Z(\rdata_LSU [1] ) );
BUF_X1 \myminixbar/_1230_ ( .A(\myminixbar/_0391_ ), .Z(\rdata_LSU [2] ) );
BUF_X1 \myminixbar/_1231_ ( .A(\myminixbar/_0394_ ), .Z(\rdata_LSU [3] ) );
BUF_X1 \myminixbar/_1232_ ( .A(\myminixbar/_0395_ ), .Z(\rdata_LSU [4] ) );
BUF_X1 \myminixbar/_1233_ ( .A(\myminixbar/_0396_ ), .Z(\rdata_LSU [5] ) );
BUF_X1 \myminixbar/_1234_ ( .A(\myminixbar/_0397_ ), .Z(\rdata_LSU [6] ) );
BUF_X1 \myminixbar/_1235_ ( .A(\myminixbar/_0398_ ), .Z(\rdata_LSU [7] ) );
BUF_X1 \myminixbar/_1236_ ( .A(\myminixbar/_0399_ ), .Z(\rdata_LSU [8] ) );
BUF_X1 \myminixbar/_1237_ ( .A(\myminixbar/_0400_ ), .Z(\rdata_LSU [9] ) );
BUF_X1 \myminixbar/_1238_ ( .A(\myminixbar/_0370_ ), .Z(\rdata_LSU [10] ) );
BUF_X1 \myminixbar/_1239_ ( .A(\myminixbar/_0371_ ), .Z(\rdata_LSU [11] ) );
BUF_X1 \myminixbar/_1240_ ( .A(\myminixbar/_0372_ ), .Z(\rdata_LSU [12] ) );
BUF_X1 \myminixbar/_1241_ ( .A(\myminixbar/_0373_ ), .Z(\rdata_LSU [13] ) );
BUF_X1 \myminixbar/_1242_ ( .A(\myminixbar/_0374_ ), .Z(\rdata_LSU [14] ) );
BUF_X1 \myminixbar/_1243_ ( .A(\myminixbar/_0375_ ), .Z(\rdata_LSU [15] ) );
BUF_X1 \myminixbar/_1244_ ( .A(\myminixbar/_0376_ ), .Z(\rdata_LSU [16] ) );
BUF_X1 \myminixbar/_1245_ ( .A(\myminixbar/_0377_ ), .Z(\rdata_LSU [17] ) );
BUF_X1 \myminixbar/_1246_ ( .A(\myminixbar/_0378_ ), .Z(\rdata_LSU [18] ) );
BUF_X1 \myminixbar/_1247_ ( .A(\myminixbar/_0379_ ), .Z(\rdata_LSU [19] ) );
BUF_X1 \myminixbar/_1248_ ( .A(\myminixbar/_0381_ ), .Z(\rdata_LSU [20] ) );
BUF_X1 \myminixbar/_1249_ ( .A(\myminixbar/_0382_ ), .Z(\rdata_LSU [21] ) );
BUF_X1 \myminixbar/_1250_ ( .A(\myminixbar/_0383_ ), .Z(\rdata_LSU [22] ) );
BUF_X1 \myminixbar/_1251_ ( .A(\myminixbar/_0384_ ), .Z(\rdata_LSU [23] ) );
BUF_X1 \myminixbar/_1252_ ( .A(\myminixbar/_0385_ ), .Z(\rdata_LSU [24] ) );
BUF_X1 \myminixbar/_1253_ ( .A(\myminixbar/_0386_ ), .Z(\rdata_LSU [25] ) );
BUF_X1 \myminixbar/_1254_ ( .A(\myminixbar/_0387_ ), .Z(\rdata_LSU [26] ) );
BUF_X1 \myminixbar/_1255_ ( .A(\myminixbar/_0388_ ), .Z(\rdata_LSU [27] ) );
BUF_X1 \myminixbar/_1256_ ( .A(\myminixbar/_0389_ ), .Z(\rdata_LSU [28] ) );
BUF_X1 \myminixbar/_1257_ ( .A(\myminixbar/_0390_ ), .Z(\rdata_LSU [29] ) );
BUF_X1 \myminixbar/_1258_ ( .A(\myminixbar/_0392_ ), .Z(\rdata_LSU [30] ) );
BUF_X1 \myminixbar/_1259_ ( .A(\myminixbar/_0393_ ), .Z(\rdata_LSU [31] ) );
BUF_X1 \myminixbar/_1260_ ( .A(\rresp_clint [0] ), .Z(\myminixbar/_0495_ ) );
BUF_X1 \myminixbar/_1261_ ( .A(\io_master_rresp [0] ), .Z(\myminixbar/_0497_ ) );
BUF_X1 \myminixbar/_1262_ ( .A(\myminixbar/_0491_ ), .Z(\rresp_IFU [0] ) );
BUF_X1 \myminixbar/_1263_ ( .A(\rresp_clint [1] ), .Z(\myminixbar/_0496_ ) );
BUF_X1 \myminixbar/_1264_ ( .A(\io_master_rresp [1] ), .Z(\myminixbar/_0498_ ) );
BUF_X1 \myminixbar/_1265_ ( .A(\myminixbar/_0492_ ), .Z(\rresp_IFU [1] ) );
BUF_X1 \myminixbar/_1266_ ( .A(\myminixbar/_0493_ ), .Z(\rresp_LSU [0] ) );
BUF_X1 \myminixbar/_1267_ ( .A(\myminixbar/_0494_ ), .Z(\rresp_LSU [1] ) );
BUF_X1 \myminixbar/_1268_ ( .A(\myminixbar/_0490_ ), .Z(io_master_rready ) );
BUF_X1 \myminixbar/_1269_ ( .A(\rid_clint [0] ), .Z(\myminixbar/_0473_ ) );
BUF_X1 \myminixbar/_1270_ ( .A(\io_master_rid [0] ), .Z(\myminixbar/_0477_ ) );
BUF_X1 \myminixbar/_1271_ ( .A(\myminixbar/_0465_ ), .Z(\rid_IFU [0] ) );
BUF_X1 \myminixbar/_1272_ ( .A(\rid_clint [1] ), .Z(\myminixbar/_0474_ ) );
BUF_X1 \myminixbar/_1273_ ( .A(\io_master_rid [1] ), .Z(\myminixbar/_0478_ ) );
BUF_X1 \myminixbar/_1274_ ( .A(\myminixbar/_0466_ ), .Z(\rid_IFU [1] ) );
BUF_X1 \myminixbar/_1275_ ( .A(\rid_clint [2] ), .Z(\myminixbar/_0475_ ) );
BUF_X1 \myminixbar/_1276_ ( .A(\io_master_rid [2] ), .Z(\myminixbar/_0479_ ) );
BUF_X1 \myminixbar/_1277_ ( .A(\myminixbar/_0467_ ), .Z(\rid_IFU [2] ) );
BUF_X1 \myminixbar/_1278_ ( .A(\rid_clint [3] ), .Z(\myminixbar/_0476_ ) );
BUF_X1 \myminixbar/_1279_ ( .A(\io_master_rid [3] ), .Z(\myminixbar/_0480_ ) );
BUF_X1 \myminixbar/_1280_ ( .A(\myminixbar/_0468_ ), .Z(\rid_IFU [3] ) );
BUF_X1 \myminixbar/_1281_ ( .A(\myminixbar/_0469_ ), .Z(\rid_LSU [0] ) );
BUF_X1 \myminixbar/_1282_ ( .A(\myminixbar/_0470_ ), .Z(\rid_LSU [1] ) );
BUF_X1 \myminixbar/_1283_ ( .A(\myminixbar/_0471_ ), .Z(\rid_LSU [2] ) );
BUF_X1 \myminixbar/_1284_ ( .A(\myminixbar/_0472_ ), .Z(\rid_LSU [3] ) );
OR2_X1 \myreg/_3474_ ( .A1(fanout_net_29 ), .A2(\myreg/_0160_ ), .ZN(\myreg/_1024_ ) );
INV_X2 \myreg/_3475_ ( .A(fanout_net_29 ), .ZN(\myreg/_1025_ ) );
BUF_X4 \myreg/_3476_ ( .A(\myreg/_1025_ ), .Z(\myreg/_1026_ ) );
BUF_X4 \myreg/_3477_ ( .A(\myreg/_1026_ ), .Z(\myreg/_1027_ ) );
OAI211_X2 \myreg/_3478_ ( .A(\myreg/_1024_ ), .B(fanout_net_38 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0192_ ), .ZN(\myreg/_1028_ ) );
INV_X1 \myreg/_3479_ ( .A(\myreg/_0128_ ), .ZN(\myreg/_1029_ ) );
AOI21_X1 \myreg/_3480_ ( .A(fanout_net_38 ), .B1(\myreg/_1029_ ), .B2(fanout_net_29 ), .ZN(\myreg/_1030_ ) );
OAI21_X1 \myreg/_3481_ ( .A(\myreg/_1030_ ), .B1(fanout_net_29 ), .B2(\myreg/_0096_ ), .ZN(\myreg/_1031_ ) );
NAND3_X1 \myreg/_3482_ ( .A1(\myreg/_1028_ ), .A2(\myreg/_1031_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1032_ ) );
OR2_X1 \myreg/_3483_ ( .A1(fanout_net_29 ), .A2(\myreg/_0032_ ), .ZN(\myreg/_1033_ ) );
OAI211_X2 \myreg/_3484_ ( .A(\myreg/_1033_ ), .B(fanout_net_38 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0064_ ), .ZN(\myreg/_1034_ ) );
INV_X1 \myreg/_3485_ ( .A(\myreg/_0480_ ), .ZN(\myreg/_1035_ ) );
AOI21_X1 \myreg/_3486_ ( .A(fanout_net_38 ), .B1(\myreg/_1035_ ), .B2(fanout_net_29 ), .ZN(\myreg/_1036_ ) );
OAI21_X1 \myreg/_3487_ ( .A(\myreg/_1036_ ), .B1(fanout_net_29 ), .B2(\myreg/_0448_ ), .ZN(\myreg/_1037_ ) );
INV_X1 \myreg/_3488_ ( .A(fanout_net_44 ), .ZN(\myreg/_1038_ ) );
BUF_X4 \myreg/_3489_ ( .A(\myreg/_1038_ ), .Z(\myreg/_1039_ ) );
BUF_X4 \myreg/_3490_ ( .A(\myreg/_1039_ ), .Z(\myreg/_1040_ ) );
NAND3_X1 \myreg/_3491_ ( .A1(\myreg/_1034_ ), .A2(\myreg/_1037_ ), .A3(\myreg/_1040_ ), .ZN(\myreg/_1041_ ) );
AND2_X1 \myreg/_3492_ ( .A1(\myreg/_1032_ ), .A2(\myreg/_1041_ ), .ZN(\myreg/_1042_ ) );
MUX2_X1 \myreg/_3493_ ( .A(\myreg/_0320_ ), .B(\myreg/_0352_ ), .S(fanout_net_29 ), .Z(\myreg/_1043_ ) );
MUX2_X1 \myreg/_3494_ ( .A(\myreg/_0384_ ), .B(\myreg/_0416_ ), .S(fanout_net_29 ), .Z(\myreg/_1044_ ) );
MUX2_X1 \myreg/_3495_ ( .A(\myreg/_1043_ ), .B(\myreg/_1044_ ), .S(fanout_net_38 ), .Z(\myreg/_1045_ ) );
MUX2_X1 \myreg/_3496_ ( .A(\myreg/_0000_ ), .B(\myreg/_0224_ ), .S(fanout_net_29 ), .Z(\myreg/_1046_ ) );
MUX2_X1 \myreg/_3497_ ( .A(\myreg/_0256_ ), .B(\myreg/_0288_ ), .S(fanout_net_29 ), .Z(\myreg/_1047_ ) );
MUX2_X1 \myreg/_3498_ ( .A(\myreg/_1046_ ), .B(\myreg/_1047_ ), .S(fanout_net_38 ), .Z(\myreg/_1048_ ) );
BUF_X4 \myreg/_3499_ ( .A(\myreg/_1039_ ), .Z(\myreg/_1049_ ) );
MUX2_X1 \myreg/_3500_ ( .A(\myreg/_1045_ ), .B(\myreg/_1048_ ), .S(\myreg/_1049_ ), .Z(\myreg/_1050_ ) );
INV_X1 \myreg/_3501_ ( .A(\myreg/_2343_ ), .ZN(\myreg/_1051_ ) );
BUF_X4 \myreg/_3502_ ( .A(\myreg/_1051_ ), .Z(\myreg/_1052_ ) );
MUX2_X1 \myreg/_3503_ ( .A(\myreg/_1042_ ), .B(\myreg/_1050_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2348_ ) );
OR2_X1 \myreg/_3504_ ( .A1(fanout_net_29 ), .A2(\myreg/_0043_ ), .ZN(\myreg/_1053_ ) );
BUF_X4 \myreg/_3505_ ( .A(\myreg/_1025_ ), .Z(\myreg/_1054_ ) );
OAI211_X2 \myreg/_3506_ ( .A(\myreg/_1053_ ), .B(fanout_net_38 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0075_ ), .ZN(\myreg/_1055_ ) );
INV_X1 \myreg/_3507_ ( .A(\myreg/_0491_ ), .ZN(\myreg/_1056_ ) );
AOI21_X1 \myreg/_3508_ ( .A(fanout_net_38 ), .B1(\myreg/_1056_ ), .B2(fanout_net_29 ), .ZN(\myreg/_1057_ ) );
OAI21_X1 \myreg/_3509_ ( .A(\myreg/_1057_ ), .B1(fanout_net_29 ), .B2(\myreg/_0459_ ), .ZN(\myreg/_1058_ ) );
AOI21_X1 \myreg/_3510_ ( .A(fanout_net_44 ), .B1(\myreg/_1055_ ), .B2(\myreg/_1058_ ), .ZN(\myreg/_1059_ ) );
OR2_X1 \myreg/_3511_ ( .A1(fanout_net_29 ), .A2(\myreg/_0171_ ), .ZN(\myreg/_1060_ ) );
OAI211_X2 \myreg/_3512_ ( .A(\myreg/_1060_ ), .B(fanout_net_38 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0203_ ), .ZN(\myreg/_1061_ ) );
INV_X1 \myreg/_3513_ ( .A(\myreg/_0139_ ), .ZN(\myreg/_1062_ ) );
AOI21_X1 \myreg/_3514_ ( .A(fanout_net_38 ), .B1(\myreg/_1062_ ), .B2(fanout_net_29 ), .ZN(\myreg/_1063_ ) );
OAI21_X1 \myreg/_3515_ ( .A(\myreg/_1063_ ), .B1(fanout_net_29 ), .B2(\myreg/_0107_ ), .ZN(\myreg/_1064_ ) );
AOI21_X1 \myreg/_3516_ ( .A(\myreg/_1039_ ), .B1(\myreg/_1061_ ), .B2(\myreg/_1064_ ), .ZN(\myreg/_1065_ ) );
OR2_X1 \myreg/_3517_ ( .A1(\myreg/_1059_ ), .A2(\myreg/_1065_ ), .ZN(\myreg/_1066_ ) );
MUX2_X1 \myreg/_3518_ ( .A(\myreg/_0331_ ), .B(\myreg/_0363_ ), .S(fanout_net_29 ), .Z(\myreg/_1067_ ) );
MUX2_X1 \myreg/_3519_ ( .A(\myreg/_0395_ ), .B(\myreg/_0427_ ), .S(fanout_net_29 ), .Z(\myreg/_1068_ ) );
MUX2_X1 \myreg/_3520_ ( .A(\myreg/_1067_ ), .B(\myreg/_1068_ ), .S(fanout_net_38 ), .Z(\myreg/_1069_ ) );
MUX2_X1 \myreg/_3521_ ( .A(\myreg/_0011_ ), .B(\myreg/_0235_ ), .S(fanout_net_29 ), .Z(\myreg/_1070_ ) );
MUX2_X1 \myreg/_3522_ ( .A(\myreg/_0267_ ), .B(\myreg/_0299_ ), .S(fanout_net_29 ), .Z(\myreg/_1071_ ) );
MUX2_X1 \myreg/_3523_ ( .A(\myreg/_1070_ ), .B(\myreg/_1071_ ), .S(fanout_net_38 ), .Z(\myreg/_1072_ ) );
MUX2_X1 \myreg/_3524_ ( .A(\myreg/_1069_ ), .B(\myreg/_1072_ ), .S(\myreg/_1049_ ), .Z(\myreg/_1073_ ) );
MUX2_X1 \myreg/_3525_ ( .A(\myreg/_1066_ ), .B(\myreg/_1073_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2359_ ) );
BUF_X2 \myreg/_3526_ ( .A(\myreg/_1025_ ), .Z(\myreg/_1074_ ) );
OR2_X1 \myreg/_3527_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0086_ ), .ZN(\myreg/_1075_ ) );
OAI211_X2 \myreg/_3528_ ( .A(\myreg/_1075_ ), .B(fanout_net_38 ), .C1(fanout_net_29 ), .C2(\myreg/_0054_ ), .ZN(\myreg/_1076_ ) );
INV_X1 \myreg/_3529_ ( .A(\myreg/_0502_ ), .ZN(\myreg/_1077_ ) );
AOI21_X1 \myreg/_3530_ ( .A(fanout_net_38 ), .B1(\myreg/_1077_ ), .B2(fanout_net_29 ), .ZN(\myreg/_1078_ ) );
OAI21_X1 \myreg/_3531_ ( .A(\myreg/_1078_ ), .B1(fanout_net_29 ), .B2(\myreg/_0470_ ), .ZN(\myreg/_1079_ ) );
NAND3_X1 \myreg/_3532_ ( .A1(\myreg/_1076_ ), .A2(\myreg/_1040_ ), .A3(\myreg/_1079_ ), .ZN(\myreg/_1080_ ) );
OR2_X1 \myreg/_3533_ ( .A1(fanout_net_29 ), .A2(\myreg/_0182_ ), .ZN(\myreg/_1081_ ) );
OAI211_X2 \myreg/_3534_ ( .A(\myreg/_1081_ ), .B(fanout_net_38 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0214_ ), .ZN(\myreg/_1082_ ) );
INV_X1 \myreg/_3535_ ( .A(\myreg/_0150_ ), .ZN(\myreg/_1083_ ) );
AOI21_X1 \myreg/_3536_ ( .A(fanout_net_38 ), .B1(\myreg/_1083_ ), .B2(fanout_net_29 ), .ZN(\myreg/_1084_ ) );
OAI21_X1 \myreg/_3537_ ( .A(\myreg/_1084_ ), .B1(fanout_net_29 ), .B2(\myreg/_0118_ ), .ZN(\myreg/_1085_ ) );
NAND3_X1 \myreg/_3538_ ( .A1(\myreg/_1082_ ), .A2(\myreg/_1085_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1086_ ) );
AND2_X1 \myreg/_3539_ ( .A1(\myreg/_1080_ ), .A2(\myreg/_1086_ ), .ZN(\myreg/_1087_ ) );
MUX2_X1 \myreg/_3540_ ( .A(\myreg/_0342_ ), .B(\myreg/_0374_ ), .S(fanout_net_29 ), .Z(\myreg/_1088_ ) );
MUX2_X1 \myreg/_3541_ ( .A(\myreg/_0406_ ), .B(\myreg/_0438_ ), .S(fanout_net_29 ), .Z(\myreg/_1089_ ) );
MUX2_X1 \myreg/_3542_ ( .A(\myreg/_1088_ ), .B(\myreg/_1089_ ), .S(fanout_net_38 ), .Z(\myreg/_1090_ ) );
MUX2_X1 \myreg/_3543_ ( .A(\myreg/_0022_ ), .B(\myreg/_0246_ ), .S(fanout_net_29 ), .Z(\myreg/_1091_ ) );
MUX2_X1 \myreg/_3544_ ( .A(\myreg/_0278_ ), .B(\myreg/_0310_ ), .S(fanout_net_30 ), .Z(\myreg/_1092_ ) );
MUX2_X1 \myreg/_3545_ ( .A(\myreg/_1091_ ), .B(\myreg/_1092_ ), .S(fanout_net_38 ), .Z(\myreg/_1093_ ) );
MUX2_X1 \myreg/_3546_ ( .A(\myreg/_1090_ ), .B(\myreg/_1093_ ), .S(\myreg/_1049_ ), .Z(\myreg/_1094_ ) );
MUX2_X1 \myreg/_3547_ ( .A(\myreg/_1087_ ), .B(\myreg/_1094_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2370_ ) );
OR2_X1 \myreg/_3548_ ( .A1(fanout_net_30 ), .A2(\myreg/_0185_ ), .ZN(\myreg/_1095_ ) );
OAI211_X2 \myreg/_3549_ ( .A(\myreg/_1095_ ), .B(fanout_net_38 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0217_ ), .ZN(\myreg/_1096_ ) );
INV_X1 \myreg/_3550_ ( .A(\myreg/_0153_ ), .ZN(\myreg/_1097_ ) );
AOI21_X1 \myreg/_3551_ ( .A(fanout_net_38 ), .B1(\myreg/_1097_ ), .B2(fanout_net_30 ), .ZN(\myreg/_1098_ ) );
OAI21_X1 \myreg/_3552_ ( .A(\myreg/_1098_ ), .B1(fanout_net_30 ), .B2(\myreg/_0121_ ), .ZN(\myreg/_1099_ ) );
NAND3_X1 \myreg/_3553_ ( .A1(\myreg/_1096_ ), .A2(\myreg/_1099_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1100_ ) );
OR2_X1 \myreg/_3554_ ( .A1(fanout_net_30 ), .A2(\myreg/_0057_ ), .ZN(\myreg/_1101_ ) );
OAI211_X2 \myreg/_3555_ ( .A(\myreg/_1101_ ), .B(fanout_net_38 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0089_ ), .ZN(\myreg/_1102_ ) );
INV_X1 \myreg/_3556_ ( .A(\myreg/_0505_ ), .ZN(\myreg/_1103_ ) );
AOI21_X1 \myreg/_3557_ ( .A(fanout_net_38 ), .B1(\myreg/_1103_ ), .B2(fanout_net_30 ), .ZN(\myreg/_1104_ ) );
OAI21_X1 \myreg/_3558_ ( .A(\myreg/_1104_ ), .B1(fanout_net_30 ), .B2(\myreg/_0473_ ), .ZN(\myreg/_1105_ ) );
NAND3_X1 \myreg/_3559_ ( .A1(\myreg/_1102_ ), .A2(\myreg/_1105_ ), .A3(\myreg/_1040_ ), .ZN(\myreg/_1106_ ) );
AND2_X1 \myreg/_3560_ ( .A1(\myreg/_1100_ ), .A2(\myreg/_1106_ ), .ZN(\myreg/_1107_ ) );
MUX2_X1 \myreg/_3561_ ( .A(\myreg/_0345_ ), .B(\myreg/_0377_ ), .S(fanout_net_30 ), .Z(\myreg/_1108_ ) );
MUX2_X1 \myreg/_3562_ ( .A(\myreg/_0409_ ), .B(\myreg/_0441_ ), .S(fanout_net_30 ), .Z(\myreg/_1109_ ) );
MUX2_X1 \myreg/_3563_ ( .A(\myreg/_1108_ ), .B(\myreg/_1109_ ), .S(fanout_net_38 ), .Z(\myreg/_1110_ ) );
MUX2_X1 \myreg/_3564_ ( .A(\myreg/_0025_ ), .B(\myreg/_0249_ ), .S(fanout_net_30 ), .Z(\myreg/_1111_ ) );
MUX2_X1 \myreg/_3565_ ( .A(\myreg/_0281_ ), .B(\myreg/_0313_ ), .S(fanout_net_30 ), .Z(\myreg/_1112_ ) );
MUX2_X1 \myreg/_3566_ ( .A(\myreg/_1111_ ), .B(\myreg/_1112_ ), .S(fanout_net_38 ), .Z(\myreg/_1113_ ) );
BUF_X4 \myreg/_3567_ ( .A(\myreg/_1039_ ), .Z(\myreg/_1114_ ) );
MUX2_X1 \myreg/_3568_ ( .A(\myreg/_1110_ ), .B(\myreg/_1113_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1115_ ) );
MUX2_X1 \myreg/_3569_ ( .A(\myreg/_1107_ ), .B(\myreg/_1115_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2373_ ) );
OR2_X1 \myreg/_3570_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0218_ ), .ZN(\myreg/_1116_ ) );
OAI211_X2 \myreg/_3571_ ( .A(\myreg/_1116_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg/_0186_ ), .ZN(\myreg/_1117_ ) );
INV_X1 \myreg/_3572_ ( .A(\myreg/_0154_ ), .ZN(\myreg/_1118_ ) );
AOI21_X1 \myreg/_3573_ ( .A(fanout_net_38 ), .B1(\myreg/_1118_ ), .B2(fanout_net_30 ), .ZN(\myreg/_1119_ ) );
OAI21_X1 \myreg/_3574_ ( .A(\myreg/_1119_ ), .B1(fanout_net_30 ), .B2(\myreg/_0122_ ), .ZN(\myreg/_1120_ ) );
NAND3_X1 \myreg/_3575_ ( .A1(\myreg/_1117_ ), .A2(fanout_net_44 ), .A3(\myreg/_1120_ ), .ZN(\myreg/_1121_ ) );
OR2_X1 \myreg/_3576_ ( .A1(fanout_net_30 ), .A2(\myreg/_0058_ ), .ZN(\myreg/_1122_ ) );
OAI211_X2 \myreg/_3577_ ( .A(\myreg/_1122_ ), .B(fanout_net_38 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0090_ ), .ZN(\myreg/_1123_ ) );
INV_X1 \myreg/_3578_ ( .A(\myreg/_0506_ ), .ZN(\myreg/_1124_ ) );
AOI21_X1 \myreg/_3579_ ( .A(fanout_net_38 ), .B1(\myreg/_1124_ ), .B2(fanout_net_30 ), .ZN(\myreg/_1125_ ) );
OAI21_X1 \myreg/_3580_ ( .A(\myreg/_1125_ ), .B1(fanout_net_30 ), .B2(\myreg/_0474_ ), .ZN(\myreg/_1126_ ) );
NAND3_X1 \myreg/_3581_ ( .A1(\myreg/_1123_ ), .A2(\myreg/_1126_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1127_ ) );
AND2_X1 \myreg/_3582_ ( .A1(\myreg/_1121_ ), .A2(\myreg/_1127_ ), .ZN(\myreg/_1128_ ) );
MUX2_X1 \myreg/_3583_ ( .A(\myreg/_0346_ ), .B(\myreg/_0378_ ), .S(fanout_net_30 ), .Z(\myreg/_1129_ ) );
MUX2_X1 \myreg/_3584_ ( .A(\myreg/_0410_ ), .B(\myreg/_0442_ ), .S(fanout_net_30 ), .Z(\myreg/_1130_ ) );
MUX2_X1 \myreg/_3585_ ( .A(\myreg/_1129_ ), .B(\myreg/_1130_ ), .S(fanout_net_38 ), .Z(\myreg/_1131_ ) );
MUX2_X1 \myreg/_3586_ ( .A(\myreg/_0026_ ), .B(\myreg/_0250_ ), .S(fanout_net_30 ), .Z(\myreg/_1132_ ) );
MUX2_X1 \myreg/_3587_ ( .A(\myreg/_0282_ ), .B(\myreg/_0314_ ), .S(fanout_net_30 ), .Z(\myreg/_1133_ ) );
MUX2_X1 \myreg/_3588_ ( .A(\myreg/_1132_ ), .B(\myreg/_1133_ ), .S(fanout_net_38 ), .Z(\myreg/_1134_ ) );
MUX2_X1 \myreg/_3589_ ( .A(\myreg/_1131_ ), .B(\myreg/_1134_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1135_ ) );
MUX2_X1 \myreg/_3590_ ( .A(\myreg/_1128_ ), .B(\myreg/_1135_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2374_ ) );
MUX2_X1 \myreg/_3591_ ( .A(\myreg/_0123_ ), .B(\myreg/_0155_ ), .S(fanout_net_30 ), .Z(\myreg/_1136_ ) );
MUX2_X1 \myreg/_3592_ ( .A(\myreg/_0187_ ), .B(\myreg/_0219_ ), .S(fanout_net_30 ), .Z(\myreg/_1137_ ) );
MUX2_X1 \myreg/_3593_ ( .A(\myreg/_1136_ ), .B(\myreg/_1137_ ), .S(fanout_net_39 ), .Z(\myreg/_1138_ ) );
MUX2_X1 \myreg/_3594_ ( .A(\myreg/_0475_ ), .B(\myreg/_0507_ ), .S(fanout_net_30 ), .Z(\myreg/_1139_ ) );
MUX2_X1 \myreg/_3595_ ( .A(\myreg/_0059_ ), .B(\myreg/_0091_ ), .S(fanout_net_30 ), .Z(\myreg/_1140_ ) );
MUX2_X1 \myreg/_3596_ ( .A(\myreg/_1139_ ), .B(\myreg/_1140_ ), .S(fanout_net_39 ), .Z(\myreg/_1141_ ) );
BUF_X4 \myreg/_3597_ ( .A(\myreg/_1038_ ), .Z(\myreg/_1142_ ) );
MUX2_X1 \myreg/_3598_ ( .A(\myreg/_1138_ ), .B(\myreg/_1141_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1143_ ) );
MUX2_X1 \myreg/_3599_ ( .A(\myreg/_0027_ ), .B(\myreg/_0283_ ), .S(fanout_net_39 ), .Z(\myreg/_1144_ ) );
MUX2_X1 \myreg/_3600_ ( .A(\myreg/_0251_ ), .B(\myreg/_0315_ ), .S(fanout_net_39 ), .Z(\myreg/_1145_ ) );
MUX2_X1 \myreg/_3601_ ( .A(\myreg/_1144_ ), .B(\myreg/_1145_ ), .S(fanout_net_30 ), .Z(\myreg/_1146_ ) );
MUX2_X1 \myreg/_3602_ ( .A(\myreg/_0347_ ), .B(\myreg/_0411_ ), .S(fanout_net_39 ), .Z(\myreg/_1147_ ) );
MUX2_X1 \myreg/_3603_ ( .A(\myreg/_0379_ ), .B(\myreg/_0443_ ), .S(fanout_net_39 ), .Z(\myreg/_1148_ ) );
MUX2_X1 \myreg/_3604_ ( .A(\myreg/_1147_ ), .B(\myreg/_1148_ ), .S(fanout_net_30 ), .Z(\myreg/_1149_ ) );
MUX2_X1 \myreg/_3605_ ( .A(\myreg/_1146_ ), .B(\myreg/_1149_ ), .S(fanout_net_44 ), .Z(\myreg/_1150_ ) );
MUX2_X1 \myreg/_3606_ ( .A(\myreg/_1143_ ), .B(\myreg/_1150_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2375_ ) );
MUX2_X1 \myreg/_3607_ ( .A(\myreg/_0124_ ), .B(\myreg/_0156_ ), .S(fanout_net_30 ), .Z(\myreg/_1151_ ) );
MUX2_X1 \myreg/_3608_ ( .A(\myreg/_0188_ ), .B(\myreg/_0220_ ), .S(fanout_net_30 ), .Z(\myreg/_1152_ ) );
MUX2_X1 \myreg/_3609_ ( .A(\myreg/_1151_ ), .B(\myreg/_1152_ ), .S(fanout_net_39 ), .Z(\myreg/_1153_ ) );
MUX2_X1 \myreg/_3610_ ( .A(\myreg/_0476_ ), .B(\myreg/_0508_ ), .S(fanout_net_30 ), .Z(\myreg/_1154_ ) );
MUX2_X1 \myreg/_3611_ ( .A(\myreg/_0060_ ), .B(\myreg/_0092_ ), .S(fanout_net_31 ), .Z(\myreg/_1155_ ) );
MUX2_X1 \myreg/_3612_ ( .A(\myreg/_1154_ ), .B(\myreg/_1155_ ), .S(fanout_net_39 ), .Z(\myreg/_1156_ ) );
MUX2_X1 \myreg/_3613_ ( .A(\myreg/_1153_ ), .B(\myreg/_1156_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1157_ ) );
MUX2_X1 \myreg/_3614_ ( .A(\myreg/_0028_ ), .B(\myreg/_0284_ ), .S(fanout_net_39 ), .Z(\myreg/_1158_ ) );
MUX2_X1 \myreg/_3615_ ( .A(\myreg/_0252_ ), .B(\myreg/_0316_ ), .S(fanout_net_39 ), .Z(\myreg/_1159_ ) );
MUX2_X1 \myreg/_3616_ ( .A(\myreg/_1158_ ), .B(\myreg/_1159_ ), .S(fanout_net_31 ), .Z(\myreg/_1160_ ) );
MUX2_X1 \myreg/_3617_ ( .A(\myreg/_0348_ ), .B(\myreg/_0412_ ), .S(fanout_net_39 ), .Z(\myreg/_1161_ ) );
MUX2_X1 \myreg/_3618_ ( .A(\myreg/_0380_ ), .B(\myreg/_0444_ ), .S(fanout_net_39 ), .Z(\myreg/_1162_ ) );
MUX2_X1 \myreg/_3619_ ( .A(\myreg/_1161_ ), .B(\myreg/_1162_ ), .S(fanout_net_31 ), .Z(\myreg/_1163_ ) );
MUX2_X1 \myreg/_3620_ ( .A(\myreg/_1160_ ), .B(\myreg/_1163_ ), .S(fanout_net_44 ), .Z(\myreg/_1164_ ) );
MUX2_X1 \myreg/_3621_ ( .A(\myreg/_1157_ ), .B(\myreg/_1164_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2376_ ) );
MUX2_X1 \myreg/_3622_ ( .A(\myreg/_0125_ ), .B(\myreg/_0157_ ), .S(fanout_net_31 ), .Z(\myreg/_1165_ ) );
MUX2_X1 \myreg/_3623_ ( .A(\myreg/_0189_ ), .B(\myreg/_0221_ ), .S(fanout_net_31 ), .Z(\myreg/_1166_ ) );
MUX2_X1 \myreg/_3624_ ( .A(\myreg/_1165_ ), .B(\myreg/_1166_ ), .S(fanout_net_39 ), .Z(\myreg/_1167_ ) );
MUX2_X1 \myreg/_3625_ ( .A(\myreg/_0477_ ), .B(\myreg/_0509_ ), .S(fanout_net_31 ), .Z(\myreg/_1168_ ) );
MUX2_X1 \myreg/_3626_ ( .A(\myreg/_0061_ ), .B(\myreg/_0093_ ), .S(fanout_net_31 ), .Z(\myreg/_1169_ ) );
MUX2_X1 \myreg/_3627_ ( .A(\myreg/_1168_ ), .B(\myreg/_1169_ ), .S(fanout_net_39 ), .Z(\myreg/_1170_ ) );
MUX2_X1 \myreg/_3628_ ( .A(\myreg/_1167_ ), .B(\myreg/_1170_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1171_ ) );
MUX2_X1 \myreg/_3629_ ( .A(\myreg/_0029_ ), .B(\myreg/_0285_ ), .S(fanout_net_39 ), .Z(\myreg/_1172_ ) );
MUX2_X1 \myreg/_3630_ ( .A(\myreg/_0253_ ), .B(\myreg/_0317_ ), .S(fanout_net_39 ), .Z(\myreg/_1173_ ) );
MUX2_X1 \myreg/_3631_ ( .A(\myreg/_1172_ ), .B(\myreg/_1173_ ), .S(fanout_net_31 ), .Z(\myreg/_1174_ ) );
MUX2_X1 \myreg/_3632_ ( .A(\myreg/_0349_ ), .B(\myreg/_0413_ ), .S(fanout_net_39 ), .Z(\myreg/_1175_ ) );
MUX2_X1 \myreg/_3633_ ( .A(\myreg/_0381_ ), .B(\myreg/_0445_ ), .S(fanout_net_39 ), .Z(\myreg/_1176_ ) );
MUX2_X1 \myreg/_3634_ ( .A(\myreg/_1175_ ), .B(\myreg/_1176_ ), .S(fanout_net_31 ), .Z(\myreg/_1177_ ) );
MUX2_X1 \myreg/_3635_ ( .A(\myreg/_1174_ ), .B(\myreg/_1177_ ), .S(fanout_net_44 ), .Z(\myreg/_1178_ ) );
MUX2_X1 \myreg/_3636_ ( .A(\myreg/_1171_ ), .B(\myreg/_1178_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2377_ ) );
OR2_X1 \myreg/_3637_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0222_ ), .ZN(\myreg/_1179_ ) );
OAI211_X2 \myreg/_3638_ ( .A(\myreg/_1179_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg/_0190_ ), .ZN(\myreg/_1180_ ) );
INV_X1 \myreg/_3639_ ( .A(\myreg/_0158_ ), .ZN(\myreg/_1181_ ) );
AOI21_X1 \myreg/_3640_ ( .A(fanout_net_39 ), .B1(\myreg/_1181_ ), .B2(fanout_net_31 ), .ZN(\myreg/_1182_ ) );
OAI21_X1 \myreg/_3641_ ( .A(\myreg/_1182_ ), .B1(fanout_net_31 ), .B2(\myreg/_0126_ ), .ZN(\myreg/_1183_ ) );
NAND3_X1 \myreg/_3642_ ( .A1(\myreg/_1180_ ), .A2(fanout_net_44 ), .A3(\myreg/_1183_ ), .ZN(\myreg/_1184_ ) );
OR2_X1 \myreg/_3643_ ( .A1(fanout_net_31 ), .A2(\myreg/_0062_ ), .ZN(\myreg/_1185_ ) );
OAI211_X2 \myreg/_3644_ ( .A(\myreg/_1185_ ), .B(fanout_net_39 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0094_ ), .ZN(\myreg/_1186_ ) );
INV_X1 \myreg/_3645_ ( .A(\myreg/_0510_ ), .ZN(\myreg/_1187_ ) );
AOI21_X1 \myreg/_3646_ ( .A(fanout_net_39 ), .B1(\myreg/_1187_ ), .B2(fanout_net_31 ), .ZN(\myreg/_1188_ ) );
OAI21_X1 \myreg/_3647_ ( .A(\myreg/_1188_ ), .B1(fanout_net_31 ), .B2(\myreg/_0478_ ), .ZN(\myreg/_1189_ ) );
NAND3_X1 \myreg/_3648_ ( .A1(\myreg/_1186_ ), .A2(\myreg/_1189_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1190_ ) );
AND2_X1 \myreg/_3649_ ( .A1(\myreg/_1184_ ), .A2(\myreg/_1190_ ), .ZN(\myreg/_1191_ ) );
MUX2_X1 \myreg/_3650_ ( .A(\myreg/_0350_ ), .B(\myreg/_0382_ ), .S(fanout_net_31 ), .Z(\myreg/_1192_ ) );
MUX2_X1 \myreg/_3651_ ( .A(\myreg/_0414_ ), .B(\myreg/_0446_ ), .S(fanout_net_31 ), .Z(\myreg/_1193_ ) );
MUX2_X1 \myreg/_3652_ ( .A(\myreg/_1192_ ), .B(\myreg/_1193_ ), .S(fanout_net_39 ), .Z(\myreg/_1194_ ) );
MUX2_X1 \myreg/_3653_ ( .A(\myreg/_0030_ ), .B(\myreg/_0254_ ), .S(fanout_net_31 ), .Z(\myreg/_1195_ ) );
MUX2_X1 \myreg/_3654_ ( .A(\myreg/_0286_ ), .B(\myreg/_0318_ ), .S(fanout_net_31 ), .Z(\myreg/_1196_ ) );
MUX2_X1 \myreg/_3655_ ( .A(\myreg/_1195_ ), .B(\myreg/_1196_ ), .S(fanout_net_39 ), .Z(\myreg/_1197_ ) );
MUX2_X1 \myreg/_3656_ ( .A(\myreg/_1194_ ), .B(\myreg/_1197_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1198_ ) );
MUX2_X1 \myreg/_3657_ ( .A(\myreg/_1191_ ), .B(\myreg/_1198_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2378_ ) );
CLKBUF_X2 \myreg/_3658_ ( .A(\myreg/_1025_ ), .Z(\myreg/_1199_ ) );
OR2_X1 \myreg/_3659_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0095_ ), .ZN(\myreg/_1200_ ) );
OAI211_X2 \myreg/_3660_ ( .A(\myreg/_1200_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg/_0063_ ), .ZN(\myreg/_1201_ ) );
INV_X1 \myreg/_3661_ ( .A(\myreg/_0511_ ), .ZN(\myreg/_1202_ ) );
AOI21_X1 \myreg/_3662_ ( .A(fanout_net_39 ), .B1(\myreg/_1202_ ), .B2(fanout_net_31 ), .ZN(\myreg/_1203_ ) );
OAI21_X1 \myreg/_3663_ ( .A(\myreg/_1203_ ), .B1(fanout_net_31 ), .B2(\myreg/_0479_ ), .ZN(\myreg/_1204_ ) );
AOI21_X1 \myreg/_3664_ ( .A(fanout_net_44 ), .B1(\myreg/_1201_ ), .B2(\myreg/_1204_ ), .ZN(\myreg/_1205_ ) );
OR2_X1 \myreg/_3665_ ( .A1(fanout_net_31 ), .A2(\myreg/_0191_ ), .ZN(\myreg/_1206_ ) );
OAI211_X2 \myreg/_3666_ ( .A(\myreg/_1206_ ), .B(fanout_net_39 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0223_ ), .ZN(\myreg/_1207_ ) );
INV_X1 \myreg/_3667_ ( .A(\myreg/_0159_ ), .ZN(\myreg/_1208_ ) );
AOI21_X1 \myreg/_3668_ ( .A(fanout_net_39 ), .B1(\myreg/_1208_ ), .B2(fanout_net_31 ), .ZN(\myreg/_1209_ ) );
OAI21_X1 \myreg/_3669_ ( .A(\myreg/_1209_ ), .B1(fanout_net_31 ), .B2(\myreg/_0127_ ), .ZN(\myreg/_1210_ ) );
AOI21_X1 \myreg/_3670_ ( .A(\myreg/_1039_ ), .B1(\myreg/_1207_ ), .B2(\myreg/_1210_ ), .ZN(\myreg/_1211_ ) );
OR2_X1 \myreg/_3671_ ( .A1(\myreg/_1205_ ), .A2(\myreg/_1211_ ), .ZN(\myreg/_1212_ ) );
MUX2_X1 \myreg/_3672_ ( .A(\myreg/_0351_ ), .B(\myreg/_0383_ ), .S(fanout_net_31 ), .Z(\myreg/_1213_ ) );
MUX2_X1 \myreg/_3673_ ( .A(\myreg/_0415_ ), .B(\myreg/_0447_ ), .S(fanout_net_31 ), .Z(\myreg/_1214_ ) );
MUX2_X1 \myreg/_3674_ ( .A(\myreg/_1213_ ), .B(\myreg/_1214_ ), .S(fanout_net_39 ), .Z(\myreg/_1215_ ) );
MUX2_X1 \myreg/_3675_ ( .A(\myreg/_0031_ ), .B(\myreg/_0255_ ), .S(fanout_net_31 ), .Z(\myreg/_1216_ ) );
MUX2_X1 \myreg/_3676_ ( .A(\myreg/_0287_ ), .B(\myreg/_0319_ ), .S(fanout_net_31 ), .Z(\myreg/_1217_ ) );
MUX2_X1 \myreg/_3677_ ( .A(\myreg/_1216_ ), .B(\myreg/_1217_ ), .S(fanout_net_39 ), .Z(\myreg/_1218_ ) );
MUX2_X1 \myreg/_3678_ ( .A(\myreg/_1215_ ), .B(\myreg/_1218_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1219_ ) );
MUX2_X1 \myreg/_3679_ ( .A(\myreg/_1212_ ), .B(\myreg/_1219_ ), .S(\myreg/_1052_ ), .Z(\myreg/_2379_ ) );
OR2_X1 \myreg/_3680_ ( .A1(fanout_net_31 ), .A2(\myreg/_0161_ ), .ZN(\myreg/_1220_ ) );
OAI211_X2 \myreg/_3681_ ( .A(\myreg/_1220_ ), .B(fanout_net_40 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0193_ ), .ZN(\myreg/_1221_ ) );
INV_X1 \myreg/_3682_ ( .A(\myreg/_0129_ ), .ZN(\myreg/_1222_ ) );
AOI21_X1 \myreg/_3683_ ( .A(fanout_net_40 ), .B1(\myreg/_1222_ ), .B2(fanout_net_32 ), .ZN(\myreg/_1223_ ) );
OAI21_X1 \myreg/_3684_ ( .A(\myreg/_1223_ ), .B1(fanout_net_32 ), .B2(\myreg/_0097_ ), .ZN(\myreg/_1224_ ) );
NAND3_X1 \myreg/_3685_ ( .A1(\myreg/_1221_ ), .A2(\myreg/_1224_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1225_ ) );
OR2_X1 \myreg/_3686_ ( .A1(fanout_net_32 ), .A2(\myreg/_0033_ ), .ZN(\myreg/_1226_ ) );
BUF_X4 \myreg/_3687_ ( .A(\myreg/_1074_ ), .Z(\myreg/_1227_ ) );
OAI211_X2 \myreg/_3688_ ( .A(\myreg/_1226_ ), .B(fanout_net_40 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0065_ ), .ZN(\myreg/_1228_ ) );
INV_X1 \myreg/_3689_ ( .A(\myreg/_0481_ ), .ZN(\myreg/_1229_ ) );
AOI21_X1 \myreg/_3690_ ( .A(fanout_net_40 ), .B1(\myreg/_1229_ ), .B2(fanout_net_32 ), .ZN(\myreg/_1230_ ) );
OAI21_X1 \myreg/_3691_ ( .A(\myreg/_1230_ ), .B1(fanout_net_32 ), .B2(\myreg/_0449_ ), .ZN(\myreg/_1231_ ) );
NAND3_X1 \myreg/_3692_ ( .A1(\myreg/_1228_ ), .A2(\myreg/_1231_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1232_ ) );
AND2_X1 \myreg/_3693_ ( .A1(\myreg/_1225_ ), .A2(\myreg/_1232_ ), .ZN(\myreg/_1233_ ) );
MUX2_X1 \myreg/_3694_ ( .A(\myreg/_0321_ ), .B(\myreg/_0353_ ), .S(fanout_net_32 ), .Z(\myreg/_1234_ ) );
MUX2_X1 \myreg/_3695_ ( .A(\myreg/_0385_ ), .B(\myreg/_0417_ ), .S(fanout_net_32 ), .Z(\myreg/_1235_ ) );
MUX2_X1 \myreg/_3696_ ( .A(\myreg/_1234_ ), .B(\myreg/_1235_ ), .S(fanout_net_40 ), .Z(\myreg/_1236_ ) );
MUX2_X1 \myreg/_3697_ ( .A(\myreg/_0001_ ), .B(\myreg/_0225_ ), .S(fanout_net_32 ), .Z(\myreg/_1237_ ) );
MUX2_X1 \myreg/_3698_ ( .A(\myreg/_0257_ ), .B(\myreg/_0289_ ), .S(fanout_net_32 ), .Z(\myreg/_1238_ ) );
MUX2_X1 \myreg/_3699_ ( .A(\myreg/_1237_ ), .B(\myreg/_1238_ ), .S(fanout_net_40 ), .Z(\myreg/_1239_ ) );
MUX2_X1 \myreg/_3700_ ( .A(\myreg/_1236_ ), .B(\myreg/_1239_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1240_ ) );
BUF_X4 \myreg/_3701_ ( .A(\myreg/_1051_ ), .Z(\myreg/_1241_ ) );
MUX2_X1 \myreg/_3702_ ( .A(\myreg/_1233_ ), .B(\myreg/_1240_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2349_ ) );
MUX2_X1 \myreg/_3703_ ( .A(\myreg/_0098_ ), .B(\myreg/_0130_ ), .S(fanout_net_32 ), .Z(\myreg/_1242_ ) );
MUX2_X1 \myreg/_3704_ ( .A(\myreg/_0162_ ), .B(\myreg/_0194_ ), .S(fanout_net_32 ), .Z(\myreg/_1243_ ) );
MUX2_X1 \myreg/_3705_ ( .A(\myreg/_1242_ ), .B(\myreg/_1243_ ), .S(fanout_net_40 ), .Z(\myreg/_1244_ ) );
MUX2_X1 \myreg/_3706_ ( .A(\myreg/_0450_ ), .B(\myreg/_0482_ ), .S(fanout_net_32 ), .Z(\myreg/_1245_ ) );
MUX2_X1 \myreg/_3707_ ( .A(\myreg/_0034_ ), .B(\myreg/_0066_ ), .S(fanout_net_32 ), .Z(\myreg/_1246_ ) );
MUX2_X1 \myreg/_3708_ ( .A(\myreg/_1245_ ), .B(\myreg/_1246_ ), .S(fanout_net_40 ), .Z(\myreg/_1247_ ) );
MUX2_X1 \myreg/_3709_ ( .A(\myreg/_1244_ ), .B(\myreg/_1247_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1248_ ) );
MUX2_X1 \myreg/_3710_ ( .A(\myreg/_0002_ ), .B(\myreg/_0258_ ), .S(fanout_net_40 ), .Z(\myreg/_1249_ ) );
MUX2_X1 \myreg/_3711_ ( .A(\myreg/_0226_ ), .B(\myreg/_0290_ ), .S(fanout_net_40 ), .Z(\myreg/_1250_ ) );
MUX2_X1 \myreg/_3712_ ( .A(\myreg/_1249_ ), .B(\myreg/_1250_ ), .S(fanout_net_32 ), .Z(\myreg/_1251_ ) );
MUX2_X1 \myreg/_3713_ ( .A(\myreg/_0322_ ), .B(\myreg/_0386_ ), .S(fanout_net_40 ), .Z(\myreg/_1252_ ) );
MUX2_X1 \myreg/_3714_ ( .A(\myreg/_0354_ ), .B(\myreg/_0418_ ), .S(fanout_net_40 ), .Z(\myreg/_1253_ ) );
MUX2_X1 \myreg/_3715_ ( .A(\myreg/_1252_ ), .B(\myreg/_1253_ ), .S(fanout_net_32 ), .Z(\myreg/_1254_ ) );
MUX2_X1 \myreg/_3716_ ( .A(\myreg/_1251_ ), .B(\myreg/_1254_ ), .S(fanout_net_44 ), .Z(\myreg/_1255_ ) );
MUX2_X1 \myreg/_3717_ ( .A(\myreg/_1248_ ), .B(\myreg/_1255_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2350_ ) );
OR2_X1 \myreg/_3718_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0067_ ), .ZN(\myreg/_1256_ ) );
OAI211_X2 \myreg/_3719_ ( .A(\myreg/_1256_ ), .B(fanout_net_40 ), .C1(fanout_net_32 ), .C2(\myreg/_0035_ ), .ZN(\myreg/_1257_ ) );
INV_X1 \myreg/_3720_ ( .A(\myreg/_0483_ ), .ZN(\myreg/_1258_ ) );
AOI21_X1 \myreg/_3721_ ( .A(fanout_net_40 ), .B1(\myreg/_1258_ ), .B2(fanout_net_32 ), .ZN(\myreg/_1259_ ) );
OAI21_X1 \myreg/_3722_ ( .A(\myreg/_1259_ ), .B1(fanout_net_32 ), .B2(\myreg/_0451_ ), .ZN(\myreg/_1260_ ) );
NAND3_X1 \myreg/_3723_ ( .A1(\myreg/_1257_ ), .A2(\myreg/_1040_ ), .A3(\myreg/_1260_ ), .ZN(\myreg/_1261_ ) );
OR2_X1 \myreg/_3724_ ( .A1(fanout_net_32 ), .A2(\myreg/_0163_ ), .ZN(\myreg/_1262_ ) );
OAI211_X2 \myreg/_3725_ ( .A(\myreg/_1262_ ), .B(fanout_net_40 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0195_ ), .ZN(\myreg/_1263_ ) );
INV_X1 \myreg/_3726_ ( .A(\myreg/_0131_ ), .ZN(\myreg/_1264_ ) );
AOI21_X1 \myreg/_3727_ ( .A(fanout_net_40 ), .B1(\myreg/_1264_ ), .B2(fanout_net_32 ), .ZN(\myreg/_1265_ ) );
OAI21_X1 \myreg/_3728_ ( .A(\myreg/_1265_ ), .B1(fanout_net_32 ), .B2(\myreg/_0099_ ), .ZN(\myreg/_1266_ ) );
NAND3_X1 \myreg/_3729_ ( .A1(\myreg/_1263_ ), .A2(\myreg/_1266_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1267_ ) );
AND2_X1 \myreg/_3730_ ( .A1(\myreg/_1261_ ), .A2(\myreg/_1267_ ), .ZN(\myreg/_1268_ ) );
MUX2_X1 \myreg/_3731_ ( .A(\myreg/_0323_ ), .B(\myreg/_0355_ ), .S(fanout_net_32 ), .Z(\myreg/_1269_ ) );
MUX2_X1 \myreg/_3732_ ( .A(\myreg/_0387_ ), .B(\myreg/_0419_ ), .S(fanout_net_32 ), .Z(\myreg/_1270_ ) );
MUX2_X1 \myreg/_3733_ ( .A(\myreg/_1269_ ), .B(\myreg/_1270_ ), .S(fanout_net_40 ), .Z(\myreg/_1271_ ) );
MUX2_X1 \myreg/_3734_ ( .A(\myreg/_0003_ ), .B(\myreg/_0227_ ), .S(fanout_net_32 ), .Z(\myreg/_1272_ ) );
MUX2_X1 \myreg/_3735_ ( .A(\myreg/_0259_ ), .B(\myreg/_0291_ ), .S(fanout_net_32 ), .Z(\myreg/_1273_ ) );
MUX2_X1 \myreg/_3736_ ( .A(\myreg/_1272_ ), .B(\myreg/_1273_ ), .S(fanout_net_40 ), .Z(\myreg/_1274_ ) );
MUX2_X1 \myreg/_3737_ ( .A(\myreg/_1271_ ), .B(\myreg/_1274_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1275_ ) );
MUX2_X1 \myreg/_3738_ ( .A(\myreg/_1268_ ), .B(\myreg/_1275_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2351_ ) );
NOR2_X1 \myreg/_3739_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0132_ ), .ZN(\myreg/_1276_ ) );
NOR2_X1 \myreg/_3740_ ( .A1(fanout_net_32 ), .A2(\myreg/_0100_ ), .ZN(\myreg/_1277_ ) );
OR3_X1 \myreg/_3741_ ( .A1(\myreg/_1276_ ), .A2(fanout_net_40 ), .A3(\myreg/_1277_ ), .ZN(\myreg/_1278_ ) );
OR2_X1 \myreg/_3742_ ( .A1(\myreg/_1025_ ), .A2(\myreg/_0196_ ), .ZN(\myreg/_1279_ ) );
OAI211_X2 \myreg/_3743_ ( .A(\myreg/_1279_ ), .B(fanout_net_40 ), .C1(fanout_net_32 ), .C2(\myreg/_0164_ ), .ZN(\myreg/_1280_ ) );
AOI21_X1 \myreg/_3744_ ( .A(\myreg/_1142_ ), .B1(\myreg/_1278_ ), .B2(\myreg/_1280_ ), .ZN(\myreg/_1281_ ) );
NOR2_X1 \myreg/_3745_ ( .A1(\myreg/_1025_ ), .A2(\myreg/_0484_ ), .ZN(\myreg/_1282_ ) );
NOR2_X1 \myreg/_3746_ ( .A1(fanout_net_32 ), .A2(\myreg/_0452_ ), .ZN(\myreg/_1283_ ) );
OR3_X1 \myreg/_3747_ ( .A1(\myreg/_1282_ ), .A2(fanout_net_40 ), .A3(\myreg/_1283_ ), .ZN(\myreg/_1284_ ) );
OR2_X1 \myreg/_3748_ ( .A1(fanout_net_32 ), .A2(\myreg/_0036_ ), .ZN(\myreg/_1285_ ) );
OAI211_X2 \myreg/_3749_ ( .A(\myreg/_1285_ ), .B(fanout_net_40 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0068_ ), .ZN(\myreg/_1286_ ) );
AOI21_X1 \myreg/_3750_ ( .A(fanout_net_44 ), .B1(\myreg/_1284_ ), .B2(\myreg/_1286_ ), .ZN(\myreg/_1287_ ) );
OR2_X1 \myreg/_3751_ ( .A1(\myreg/_1281_ ), .A2(\myreg/_1287_ ), .ZN(\myreg/_1288_ ) );
MUX2_X1 \myreg/_3752_ ( .A(\myreg/_0324_ ), .B(\myreg/_0356_ ), .S(fanout_net_32 ), .Z(\myreg/_1289_ ) );
MUX2_X1 \myreg/_3753_ ( .A(\myreg/_0388_ ), .B(\myreg/_0420_ ), .S(fanout_net_33 ), .Z(\myreg/_1290_ ) );
MUX2_X1 \myreg/_3754_ ( .A(\myreg/_1289_ ), .B(\myreg/_1290_ ), .S(fanout_net_40 ), .Z(\myreg/_1291_ ) );
MUX2_X1 \myreg/_3755_ ( .A(\myreg/_0004_ ), .B(\myreg/_0228_ ), .S(fanout_net_33 ), .Z(\myreg/_1292_ ) );
MUX2_X1 \myreg/_3756_ ( .A(\myreg/_0260_ ), .B(\myreg/_0292_ ), .S(fanout_net_33 ), .Z(\myreg/_1293_ ) );
MUX2_X1 \myreg/_3757_ ( .A(\myreg/_1292_ ), .B(\myreg/_1293_ ), .S(fanout_net_40 ), .Z(\myreg/_1294_ ) );
MUX2_X1 \myreg/_3758_ ( .A(\myreg/_1291_ ), .B(\myreg/_1294_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1295_ ) );
MUX2_X1 \myreg/_3759_ ( .A(\myreg/_1288_ ), .B(\myreg/_1295_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2352_ ) );
OR2_X1 \myreg/_3760_ ( .A1(fanout_net_33 ), .A2(\myreg/_0037_ ), .ZN(\myreg/_1296_ ) );
OAI211_X2 \myreg/_3761_ ( .A(\myreg/_1296_ ), .B(fanout_net_40 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0069_ ), .ZN(\myreg/_1297_ ) );
INV_X1 \myreg/_3762_ ( .A(\myreg/_0485_ ), .ZN(\myreg/_1298_ ) );
AOI21_X1 \myreg/_3763_ ( .A(fanout_net_40 ), .B1(\myreg/_1298_ ), .B2(fanout_net_33 ), .ZN(\myreg/_1299_ ) );
OAI21_X1 \myreg/_3764_ ( .A(\myreg/_1299_ ), .B1(fanout_net_33 ), .B2(\myreg/_0453_ ), .ZN(\myreg/_1300_ ) );
AOI21_X1 \myreg/_3765_ ( .A(fanout_net_44 ), .B1(\myreg/_1297_ ), .B2(\myreg/_1300_ ), .ZN(\myreg/_1301_ ) );
OR2_X1 \myreg/_3766_ ( .A1(fanout_net_33 ), .A2(\myreg/_0165_ ), .ZN(\myreg/_1302_ ) );
OAI211_X2 \myreg/_3767_ ( .A(\myreg/_1302_ ), .B(fanout_net_40 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0197_ ), .ZN(\myreg/_1303_ ) );
INV_X1 \myreg/_3768_ ( .A(\myreg/_0133_ ), .ZN(\myreg/_1304_ ) );
AOI21_X1 \myreg/_3769_ ( .A(fanout_net_40 ), .B1(\myreg/_1304_ ), .B2(fanout_net_33 ), .ZN(\myreg/_1305_ ) );
OAI21_X1 \myreg/_3770_ ( .A(\myreg/_1305_ ), .B1(fanout_net_33 ), .B2(\myreg/_0101_ ), .ZN(\myreg/_1306_ ) );
AOI21_X1 \myreg/_3771_ ( .A(\myreg/_1039_ ), .B1(\myreg/_1303_ ), .B2(\myreg/_1306_ ), .ZN(\myreg/_1307_ ) );
OR2_X1 \myreg/_3772_ ( .A1(\myreg/_1301_ ), .A2(\myreg/_1307_ ), .ZN(\myreg/_1308_ ) );
MUX2_X1 \myreg/_3773_ ( .A(\myreg/_0325_ ), .B(\myreg/_0357_ ), .S(fanout_net_33 ), .Z(\myreg/_1309_ ) );
MUX2_X1 \myreg/_3774_ ( .A(\myreg/_0389_ ), .B(\myreg/_0421_ ), .S(fanout_net_33 ), .Z(\myreg/_1310_ ) );
MUX2_X1 \myreg/_3775_ ( .A(\myreg/_1309_ ), .B(\myreg/_1310_ ), .S(fanout_net_40 ), .Z(\myreg/_1311_ ) );
MUX2_X1 \myreg/_3776_ ( .A(\myreg/_0005_ ), .B(\myreg/_0229_ ), .S(fanout_net_33 ), .Z(\myreg/_1312_ ) );
MUX2_X1 \myreg/_3777_ ( .A(\myreg/_0261_ ), .B(\myreg/_0293_ ), .S(fanout_net_33 ), .Z(\myreg/_1313_ ) );
MUX2_X1 \myreg/_3778_ ( .A(\myreg/_1312_ ), .B(\myreg/_1313_ ), .S(fanout_net_40 ), .Z(\myreg/_1314_ ) );
MUX2_X1 \myreg/_3779_ ( .A(\myreg/_1311_ ), .B(\myreg/_1314_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1315_ ) );
MUX2_X1 \myreg/_3780_ ( .A(\myreg/_1308_ ), .B(\myreg/_1315_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2353_ ) );
MUX2_X1 \myreg/_3781_ ( .A(\myreg/_0102_ ), .B(\myreg/_0134_ ), .S(fanout_net_33 ), .Z(\myreg/_1316_ ) );
MUX2_X1 \myreg/_3782_ ( .A(\myreg/_0166_ ), .B(\myreg/_0198_ ), .S(fanout_net_33 ), .Z(\myreg/_1317_ ) );
MUX2_X1 \myreg/_3783_ ( .A(\myreg/_1316_ ), .B(\myreg/_1317_ ), .S(fanout_net_41 ), .Z(\myreg/_1318_ ) );
MUX2_X1 \myreg/_3784_ ( .A(\myreg/_0454_ ), .B(\myreg/_0486_ ), .S(fanout_net_33 ), .Z(\myreg/_1319_ ) );
MUX2_X1 \myreg/_3785_ ( .A(\myreg/_0038_ ), .B(\myreg/_0070_ ), .S(fanout_net_33 ), .Z(\myreg/_1320_ ) );
MUX2_X1 \myreg/_3786_ ( .A(\myreg/_1319_ ), .B(\myreg/_1320_ ), .S(fanout_net_41 ), .Z(\myreg/_1321_ ) );
MUX2_X1 \myreg/_3787_ ( .A(\myreg/_1318_ ), .B(\myreg/_1321_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1322_ ) );
MUX2_X1 \myreg/_3788_ ( .A(\myreg/_0006_ ), .B(\myreg/_0262_ ), .S(fanout_net_41 ), .Z(\myreg/_1323_ ) );
MUX2_X1 \myreg/_3789_ ( .A(\myreg/_0230_ ), .B(\myreg/_0294_ ), .S(fanout_net_41 ), .Z(\myreg/_1324_ ) );
MUX2_X1 \myreg/_3790_ ( .A(\myreg/_1323_ ), .B(\myreg/_1324_ ), .S(fanout_net_33 ), .Z(\myreg/_1325_ ) );
MUX2_X1 \myreg/_3791_ ( .A(\myreg/_0326_ ), .B(\myreg/_0390_ ), .S(fanout_net_41 ), .Z(\myreg/_1326_ ) );
MUX2_X1 \myreg/_3792_ ( .A(\myreg/_0358_ ), .B(\myreg/_0422_ ), .S(fanout_net_41 ), .Z(\myreg/_1327_ ) );
MUX2_X1 \myreg/_3793_ ( .A(\myreg/_1326_ ), .B(\myreg/_1327_ ), .S(fanout_net_33 ), .Z(\myreg/_1328_ ) );
MUX2_X1 \myreg/_3794_ ( .A(\myreg/_1325_ ), .B(\myreg/_1328_ ), .S(fanout_net_44 ), .Z(\myreg/_1329_ ) );
MUX2_X1 \myreg/_3795_ ( .A(\myreg/_1322_ ), .B(\myreg/_1329_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2354_ ) );
OR2_X1 \myreg/_3796_ ( .A1(fanout_net_33 ), .A2(\myreg/_0167_ ), .ZN(\myreg/_1330_ ) );
OAI211_X2 \myreg/_3797_ ( .A(\myreg/_1330_ ), .B(fanout_net_41 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0199_ ), .ZN(\myreg/_1331_ ) );
INV_X1 \myreg/_3798_ ( .A(\myreg/_0135_ ), .ZN(\myreg/_1332_ ) );
AOI21_X1 \myreg/_3799_ ( .A(fanout_net_41 ), .B1(\myreg/_1332_ ), .B2(fanout_net_33 ), .ZN(\myreg/_1333_ ) );
OAI21_X1 \myreg/_3800_ ( .A(\myreg/_1333_ ), .B1(fanout_net_33 ), .B2(\myreg/_0103_ ), .ZN(\myreg/_1334_ ) );
NAND3_X1 \myreg/_3801_ ( .A1(\myreg/_1331_ ), .A2(\myreg/_1334_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1335_ ) );
OR2_X1 \myreg/_3802_ ( .A1(fanout_net_33 ), .A2(\myreg/_0039_ ), .ZN(\myreg/_1336_ ) );
OAI211_X2 \myreg/_3803_ ( .A(\myreg/_1336_ ), .B(fanout_net_41 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0071_ ), .ZN(\myreg/_1337_ ) );
INV_X1 \myreg/_3804_ ( .A(\myreg/_0487_ ), .ZN(\myreg/_1338_ ) );
AOI21_X1 \myreg/_3805_ ( .A(fanout_net_41 ), .B1(\myreg/_1338_ ), .B2(fanout_net_33 ), .ZN(\myreg/_1339_ ) );
OAI21_X1 \myreg/_3806_ ( .A(\myreg/_1339_ ), .B1(fanout_net_33 ), .B2(\myreg/_0455_ ), .ZN(\myreg/_1340_ ) );
NAND3_X1 \myreg/_3807_ ( .A1(\myreg/_1337_ ), .A2(\myreg/_1340_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1341_ ) );
AND2_X1 \myreg/_3808_ ( .A1(\myreg/_1335_ ), .A2(\myreg/_1341_ ), .ZN(\myreg/_1342_ ) );
MUX2_X1 \myreg/_3809_ ( .A(\myreg/_0327_ ), .B(\myreg/_0359_ ), .S(fanout_net_33 ), .Z(\myreg/_1343_ ) );
MUX2_X1 \myreg/_3810_ ( .A(\myreg/_0391_ ), .B(\myreg/_0423_ ), .S(fanout_net_33 ), .Z(\myreg/_1344_ ) );
MUX2_X1 \myreg/_3811_ ( .A(\myreg/_1343_ ), .B(\myreg/_1344_ ), .S(fanout_net_41 ), .Z(\myreg/_1345_ ) );
MUX2_X1 \myreg/_3812_ ( .A(\myreg/_0007_ ), .B(\myreg/_0231_ ), .S(fanout_net_33 ), .Z(\myreg/_1346_ ) );
MUX2_X1 \myreg/_3813_ ( .A(\myreg/_0263_ ), .B(\myreg/_0295_ ), .S(fanout_net_33 ), .Z(\myreg/_1347_ ) );
MUX2_X1 \myreg/_3814_ ( .A(\myreg/_1346_ ), .B(\myreg/_1347_ ), .S(fanout_net_41 ), .Z(\myreg/_1348_ ) );
MUX2_X1 \myreg/_3815_ ( .A(\myreg/_1345_ ), .B(\myreg/_1348_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1349_ ) );
MUX2_X1 \myreg/_3816_ ( .A(\myreg/_1342_ ), .B(\myreg/_1349_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2355_ ) );
OR2_X1 \myreg/_3817_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0072_ ), .ZN(\myreg/_1350_ ) );
OAI211_X2 \myreg/_3818_ ( .A(\myreg/_1350_ ), .B(fanout_net_41 ), .C1(fanout_net_33 ), .C2(\myreg/_0040_ ), .ZN(\myreg/_1351_ ) );
INV_X1 \myreg/_3819_ ( .A(\myreg/_0488_ ), .ZN(\myreg/_1352_ ) );
AOI21_X1 \myreg/_3820_ ( .A(fanout_net_41 ), .B1(\myreg/_1352_ ), .B2(fanout_net_34 ), .ZN(\myreg/_1353_ ) );
OAI21_X1 \myreg/_3821_ ( .A(\myreg/_1353_ ), .B1(fanout_net_34 ), .B2(\myreg/_0456_ ), .ZN(\myreg/_1354_ ) );
AOI21_X1 \myreg/_3822_ ( .A(fanout_net_44 ), .B1(\myreg/_1351_ ), .B2(\myreg/_1354_ ), .ZN(\myreg/_1355_ ) );
OR2_X1 \myreg/_3823_ ( .A1(fanout_net_34 ), .A2(\myreg/_0168_ ), .ZN(\myreg/_1356_ ) );
OAI211_X2 \myreg/_3824_ ( .A(\myreg/_1356_ ), .B(fanout_net_41 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0200_ ), .ZN(\myreg/_1357_ ) );
INV_X1 \myreg/_3825_ ( .A(\myreg/_0136_ ), .ZN(\myreg/_1358_ ) );
AOI21_X1 \myreg/_3826_ ( .A(fanout_net_41 ), .B1(\myreg/_1358_ ), .B2(fanout_net_34 ), .ZN(\myreg/_1359_ ) );
OAI21_X1 \myreg/_3827_ ( .A(\myreg/_1359_ ), .B1(fanout_net_34 ), .B2(\myreg/_0104_ ), .ZN(\myreg/_1360_ ) );
AOI21_X1 \myreg/_3828_ ( .A(\myreg/_1039_ ), .B1(\myreg/_1357_ ), .B2(\myreg/_1360_ ), .ZN(\myreg/_1361_ ) );
OR2_X1 \myreg/_3829_ ( .A1(\myreg/_1355_ ), .A2(\myreg/_1361_ ), .ZN(\myreg/_1362_ ) );
MUX2_X1 \myreg/_3830_ ( .A(\myreg/_0328_ ), .B(\myreg/_0360_ ), .S(fanout_net_34 ), .Z(\myreg/_1363_ ) );
MUX2_X1 \myreg/_3831_ ( .A(\myreg/_0392_ ), .B(\myreg/_0424_ ), .S(fanout_net_34 ), .Z(\myreg/_1364_ ) );
MUX2_X1 \myreg/_3832_ ( .A(\myreg/_1363_ ), .B(\myreg/_1364_ ), .S(fanout_net_41 ), .Z(\myreg/_1365_ ) );
MUX2_X1 \myreg/_3833_ ( .A(\myreg/_0008_ ), .B(\myreg/_0232_ ), .S(fanout_net_34 ), .Z(\myreg/_1366_ ) );
MUX2_X1 \myreg/_3834_ ( .A(\myreg/_0264_ ), .B(\myreg/_0296_ ), .S(fanout_net_34 ), .Z(\myreg/_1367_ ) );
MUX2_X1 \myreg/_3835_ ( .A(\myreg/_1366_ ), .B(\myreg/_1367_ ), .S(fanout_net_41 ), .Z(\myreg/_1368_ ) );
MUX2_X1 \myreg/_3836_ ( .A(\myreg/_1365_ ), .B(\myreg/_1368_ ), .S(\myreg/_1114_ ), .Z(\myreg/_1369_ ) );
MUX2_X1 \myreg/_3837_ ( .A(\myreg/_1362_ ), .B(\myreg/_1369_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2356_ ) );
OR2_X1 \myreg/_3838_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0201_ ), .ZN(\myreg/_1370_ ) );
OAI211_X2 \myreg/_3839_ ( .A(\myreg/_1370_ ), .B(fanout_net_41 ), .C1(fanout_net_34 ), .C2(\myreg/_0169_ ), .ZN(\myreg/_1371_ ) );
INV_X1 \myreg/_3840_ ( .A(\myreg/_0137_ ), .ZN(\myreg/_1372_ ) );
AOI21_X1 \myreg/_3841_ ( .A(fanout_net_41 ), .B1(\myreg/_1372_ ), .B2(fanout_net_34 ), .ZN(\myreg/_1373_ ) );
OAI21_X1 \myreg/_3842_ ( .A(\myreg/_1373_ ), .B1(fanout_net_34 ), .B2(\myreg/_0105_ ), .ZN(\myreg/_1374_ ) );
NAND3_X1 \myreg/_3843_ ( .A1(\myreg/_1371_ ), .A2(fanout_net_44 ), .A3(\myreg/_1374_ ), .ZN(\myreg/_1375_ ) );
OR2_X1 \myreg/_3844_ ( .A1(fanout_net_34 ), .A2(\myreg/_0041_ ), .ZN(\myreg/_1376_ ) );
OAI211_X2 \myreg/_3845_ ( .A(\myreg/_1376_ ), .B(fanout_net_41 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0073_ ), .ZN(\myreg/_1377_ ) );
INV_X1 \myreg/_3846_ ( .A(\myreg/_0489_ ), .ZN(\myreg/_1378_ ) );
AOI21_X1 \myreg/_3847_ ( .A(fanout_net_41 ), .B1(\myreg/_1378_ ), .B2(fanout_net_34 ), .ZN(\myreg/_1379_ ) );
OAI21_X1 \myreg/_3848_ ( .A(\myreg/_1379_ ), .B1(fanout_net_34 ), .B2(\myreg/_0457_ ), .ZN(\myreg/_1380_ ) );
NAND3_X1 \myreg/_3849_ ( .A1(\myreg/_1377_ ), .A2(\myreg/_1380_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1381_ ) );
AND2_X1 \myreg/_3850_ ( .A1(\myreg/_1375_ ), .A2(\myreg/_1381_ ), .ZN(\myreg/_1382_ ) );
MUX2_X1 \myreg/_3851_ ( .A(\myreg/_0329_ ), .B(\myreg/_0361_ ), .S(fanout_net_34 ), .Z(\myreg/_1383_ ) );
MUX2_X1 \myreg/_3852_ ( .A(\myreg/_0393_ ), .B(\myreg/_0425_ ), .S(fanout_net_34 ), .Z(\myreg/_1384_ ) );
MUX2_X1 \myreg/_3853_ ( .A(\myreg/_1383_ ), .B(\myreg/_1384_ ), .S(fanout_net_41 ), .Z(\myreg/_1385_ ) );
MUX2_X1 \myreg/_3854_ ( .A(\myreg/_0009_ ), .B(\myreg/_0233_ ), .S(fanout_net_34 ), .Z(\myreg/_1386_ ) );
MUX2_X1 \myreg/_3855_ ( .A(\myreg/_0265_ ), .B(\myreg/_0297_ ), .S(fanout_net_34 ), .Z(\myreg/_1387_ ) );
MUX2_X1 \myreg/_3856_ ( .A(\myreg/_1386_ ), .B(\myreg/_1387_ ), .S(fanout_net_41 ), .Z(\myreg/_1388_ ) );
BUF_X4 \myreg/_3857_ ( .A(\myreg/_1039_ ), .Z(\myreg/_1389_ ) );
MUX2_X1 \myreg/_3858_ ( .A(\myreg/_1385_ ), .B(\myreg/_1388_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1390_ ) );
MUX2_X1 \myreg/_3859_ ( .A(\myreg/_1382_ ), .B(\myreg/_1390_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2357_ ) );
NOR2_X1 \myreg/_3860_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0490_ ), .ZN(\myreg/_1391_ ) );
NOR2_X1 \myreg/_3861_ ( .A1(fanout_net_34 ), .A2(\myreg/_0458_ ), .ZN(\myreg/_1392_ ) );
OR3_X1 \myreg/_3862_ ( .A1(\myreg/_1391_ ), .A2(fanout_net_41 ), .A3(\myreg/_1392_ ), .ZN(\myreg/_1393_ ) );
OR2_X1 \myreg/_3863_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0074_ ), .ZN(\myreg/_1394_ ) );
OAI211_X2 \myreg/_3864_ ( .A(\myreg/_1394_ ), .B(fanout_net_41 ), .C1(fanout_net_34 ), .C2(\myreg/_0042_ ), .ZN(\myreg/_1395_ ) );
NAND3_X1 \myreg/_3865_ ( .A1(\myreg/_1393_ ), .A2(\myreg/_1395_ ), .A3(\myreg/_1040_ ), .ZN(\myreg/_1396_ ) );
NOR2_X1 \myreg/_3866_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0138_ ), .ZN(\myreg/_1397_ ) );
NOR2_X1 \myreg/_3867_ ( .A1(fanout_net_34 ), .A2(\myreg/_0106_ ), .ZN(\myreg/_1398_ ) );
OR3_X1 \myreg/_3868_ ( .A1(\myreg/_1397_ ), .A2(fanout_net_41 ), .A3(\myreg/_1398_ ), .ZN(\myreg/_1399_ ) );
OR2_X1 \myreg/_3869_ ( .A1(fanout_net_34 ), .A2(\myreg/_0170_ ), .ZN(\myreg/_1400_ ) );
OAI211_X2 \myreg/_3870_ ( .A(\myreg/_1400_ ), .B(fanout_net_41 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0202_ ), .ZN(\myreg/_1401_ ) );
NAND3_X1 \myreg/_3871_ ( .A1(\myreg/_1399_ ), .A2(fanout_net_44 ), .A3(\myreg/_1401_ ), .ZN(\myreg/_1402_ ) );
AND2_X1 \myreg/_3872_ ( .A1(\myreg/_1396_ ), .A2(\myreg/_1402_ ), .ZN(\myreg/_1403_ ) );
MUX2_X1 \myreg/_3873_ ( .A(\myreg/_0330_ ), .B(\myreg/_0362_ ), .S(fanout_net_34 ), .Z(\myreg/_1404_ ) );
MUX2_X1 \myreg/_3874_ ( .A(\myreg/_0394_ ), .B(\myreg/_0426_ ), .S(fanout_net_34 ), .Z(\myreg/_1405_ ) );
MUX2_X1 \myreg/_3875_ ( .A(\myreg/_1404_ ), .B(\myreg/_1405_ ), .S(fanout_net_41 ), .Z(\myreg/_1406_ ) );
MUX2_X1 \myreg/_3876_ ( .A(\myreg/_0010_ ), .B(\myreg/_0234_ ), .S(fanout_net_34 ), .Z(\myreg/_1407_ ) );
MUX2_X1 \myreg/_3877_ ( .A(\myreg/_0266_ ), .B(\myreg/_0298_ ), .S(fanout_net_34 ), .Z(\myreg/_1408_ ) );
MUX2_X1 \myreg/_3878_ ( .A(\myreg/_1407_ ), .B(\myreg/_1408_ ), .S(fanout_net_41 ), .Z(\myreg/_1409_ ) );
MUX2_X1 \myreg/_3879_ ( .A(\myreg/_1406_ ), .B(\myreg/_1409_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1410_ ) );
MUX2_X1 \myreg/_3880_ ( .A(\myreg/_1403_ ), .B(\myreg/_1410_ ), .S(\myreg/_1241_ ), .Z(\myreg/_2358_ ) );
NOR2_X1 \myreg/_3881_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0140_ ), .ZN(\myreg/_1411_ ) );
NOR2_X1 \myreg/_3882_ ( .A1(fanout_net_34 ), .A2(\myreg/_0108_ ), .ZN(\myreg/_1412_ ) );
OR3_X1 \myreg/_3883_ ( .A1(\myreg/_1411_ ), .A2(fanout_net_42 ), .A3(\myreg/_1412_ ), .ZN(\myreg/_1413_ ) );
OR2_X1 \myreg/_3884_ ( .A1(fanout_net_34 ), .A2(\myreg/_0172_ ), .ZN(\myreg/_1414_ ) );
OAI211_X2 \myreg/_3885_ ( .A(\myreg/_1414_ ), .B(fanout_net_42 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0204_ ), .ZN(\myreg/_1415_ ) );
NAND3_X1 \myreg/_3886_ ( .A1(\myreg/_1413_ ), .A2(fanout_net_44 ), .A3(\myreg/_1415_ ), .ZN(\myreg/_1416_ ) );
NOR2_X1 \myreg/_3887_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0492_ ), .ZN(\myreg/_1417_ ) );
NOR2_X1 \myreg/_3888_ ( .A1(fanout_net_34 ), .A2(\myreg/_0460_ ), .ZN(\myreg/_1418_ ) );
OR3_X1 \myreg/_3889_ ( .A1(\myreg/_1417_ ), .A2(fanout_net_42 ), .A3(\myreg/_1418_ ), .ZN(\myreg/_1419_ ) );
OR2_X1 \myreg/_3890_ ( .A1(fanout_net_35 ), .A2(\myreg/_0044_ ), .ZN(\myreg/_1420_ ) );
OAI211_X2 \myreg/_3891_ ( .A(\myreg/_1420_ ), .B(fanout_net_42 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0076_ ), .ZN(\myreg/_1421_ ) );
NAND3_X1 \myreg/_3892_ ( .A1(\myreg/_1419_ ), .A2(\myreg/_1040_ ), .A3(\myreg/_1421_ ), .ZN(\myreg/_1422_ ) );
AND2_X1 \myreg/_3893_ ( .A1(\myreg/_1416_ ), .A2(\myreg/_1422_ ), .ZN(\myreg/_1423_ ) );
MUX2_X1 \myreg/_3894_ ( .A(\myreg/_0332_ ), .B(\myreg/_0364_ ), .S(fanout_net_35 ), .Z(\myreg/_1424_ ) );
MUX2_X1 \myreg/_3895_ ( .A(\myreg/_0396_ ), .B(\myreg/_0428_ ), .S(fanout_net_35 ), .Z(\myreg/_1425_ ) );
MUX2_X1 \myreg/_3896_ ( .A(\myreg/_1424_ ), .B(\myreg/_1425_ ), .S(fanout_net_42 ), .Z(\myreg/_1426_ ) );
MUX2_X1 \myreg/_3897_ ( .A(\myreg/_0012_ ), .B(\myreg/_0236_ ), .S(fanout_net_35 ), .Z(\myreg/_1427_ ) );
MUX2_X1 \myreg/_3898_ ( .A(\myreg/_0268_ ), .B(\myreg/_0300_ ), .S(fanout_net_35 ), .Z(\myreg/_1428_ ) );
MUX2_X1 \myreg/_3899_ ( .A(\myreg/_1427_ ), .B(\myreg/_1428_ ), .S(fanout_net_42 ), .Z(\myreg/_1429_ ) );
MUX2_X1 \myreg/_3900_ ( .A(\myreg/_1426_ ), .B(\myreg/_1429_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1430_ ) );
BUF_X4 \myreg/_3901_ ( .A(\myreg/_1051_ ), .Z(\myreg/_1431_ ) );
MUX2_X1 \myreg/_3902_ ( .A(\myreg/_1423_ ), .B(\myreg/_1430_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2360_ ) );
NOR2_X1 \myreg/_3903_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0493_ ), .ZN(\myreg/_1432_ ) );
NOR2_X1 \myreg/_3904_ ( .A1(fanout_net_35 ), .A2(\myreg/_0461_ ), .ZN(\myreg/_1433_ ) );
OR3_X1 \myreg/_3905_ ( .A1(\myreg/_1432_ ), .A2(fanout_net_42 ), .A3(\myreg/_1433_ ), .ZN(\myreg/_1434_ ) );
OR2_X1 \myreg/_3906_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0077_ ), .ZN(\myreg/_1435_ ) );
OAI211_X2 \myreg/_3907_ ( .A(\myreg/_1435_ ), .B(fanout_net_42 ), .C1(fanout_net_35 ), .C2(\myreg/_0045_ ), .ZN(\myreg/_1436_ ) );
NAND3_X1 \myreg/_3908_ ( .A1(\myreg/_1434_ ), .A2(\myreg/_1436_ ), .A3(\myreg/_1040_ ), .ZN(\myreg/_1437_ ) );
NOR2_X1 \myreg/_3909_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0141_ ), .ZN(\myreg/_1438_ ) );
NOR2_X1 \myreg/_3910_ ( .A1(fanout_net_35 ), .A2(\myreg/_0109_ ), .ZN(\myreg/_1439_ ) );
OR3_X1 \myreg/_3911_ ( .A1(\myreg/_1438_ ), .A2(fanout_net_42 ), .A3(\myreg/_1439_ ), .ZN(\myreg/_1440_ ) );
OR2_X1 \myreg/_3912_ ( .A1(fanout_net_35 ), .A2(\myreg/_0173_ ), .ZN(\myreg/_1441_ ) );
OAI211_X2 \myreg/_3913_ ( .A(\myreg/_1441_ ), .B(fanout_net_42 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0205_ ), .ZN(\myreg/_1442_ ) );
NAND3_X1 \myreg/_3914_ ( .A1(\myreg/_1440_ ), .A2(fanout_net_44 ), .A3(\myreg/_1442_ ), .ZN(\myreg/_1443_ ) );
AND2_X1 \myreg/_3915_ ( .A1(\myreg/_1437_ ), .A2(\myreg/_1443_ ), .ZN(\myreg/_1444_ ) );
MUX2_X1 \myreg/_3916_ ( .A(\myreg/_0333_ ), .B(\myreg/_0365_ ), .S(fanout_net_35 ), .Z(\myreg/_1445_ ) );
MUX2_X1 \myreg/_3917_ ( .A(\myreg/_0397_ ), .B(\myreg/_0429_ ), .S(fanout_net_35 ), .Z(\myreg/_1446_ ) );
MUX2_X1 \myreg/_3918_ ( .A(\myreg/_1445_ ), .B(\myreg/_1446_ ), .S(fanout_net_42 ), .Z(\myreg/_1447_ ) );
MUX2_X1 \myreg/_3919_ ( .A(\myreg/_0013_ ), .B(\myreg/_0237_ ), .S(fanout_net_35 ), .Z(\myreg/_1448_ ) );
MUX2_X1 \myreg/_3920_ ( .A(\myreg/_0269_ ), .B(\myreg/_0301_ ), .S(fanout_net_35 ), .Z(\myreg/_1449_ ) );
MUX2_X1 \myreg/_3921_ ( .A(\myreg/_1448_ ), .B(\myreg/_1449_ ), .S(fanout_net_42 ), .Z(\myreg/_1450_ ) );
MUX2_X1 \myreg/_3922_ ( .A(\myreg/_1447_ ), .B(\myreg/_1450_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1451_ ) );
MUX2_X1 \myreg/_3923_ ( .A(\myreg/_1444_ ), .B(\myreg/_1451_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2361_ ) );
OR2_X1 \myreg/_3924_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0078_ ), .ZN(\myreg/_1452_ ) );
OAI211_X2 \myreg/_3925_ ( .A(\myreg/_1452_ ), .B(fanout_net_42 ), .C1(fanout_net_35 ), .C2(\myreg/_0046_ ), .ZN(\myreg/_1453_ ) );
INV_X1 \myreg/_3926_ ( .A(\myreg/_0494_ ), .ZN(\myreg/_1454_ ) );
AOI21_X1 \myreg/_3927_ ( .A(fanout_net_42 ), .B1(\myreg/_1454_ ), .B2(fanout_net_35 ), .ZN(\myreg/_1455_ ) );
OAI21_X1 \myreg/_3928_ ( .A(\myreg/_1455_ ), .B1(fanout_net_35 ), .B2(\myreg/_0462_ ), .ZN(\myreg/_1456_ ) );
NAND3_X1 \myreg/_3929_ ( .A1(\myreg/_1453_ ), .A2(\myreg/_1040_ ), .A3(\myreg/_1456_ ), .ZN(\myreg/_1457_ ) );
OR2_X1 \myreg/_3930_ ( .A1(fanout_net_35 ), .A2(\myreg/_0174_ ), .ZN(\myreg/_1458_ ) );
OAI211_X2 \myreg/_3931_ ( .A(\myreg/_1458_ ), .B(fanout_net_42 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0206_ ), .ZN(\myreg/_1459_ ) );
INV_X1 \myreg/_3932_ ( .A(\myreg/_0142_ ), .ZN(\myreg/_1460_ ) );
AOI21_X1 \myreg/_3933_ ( .A(fanout_net_42 ), .B1(\myreg/_1460_ ), .B2(fanout_net_35 ), .ZN(\myreg/_1461_ ) );
OAI21_X1 \myreg/_3934_ ( .A(\myreg/_1461_ ), .B1(fanout_net_35 ), .B2(\myreg/_0110_ ), .ZN(\myreg/_1462_ ) );
NAND3_X1 \myreg/_3935_ ( .A1(\myreg/_1459_ ), .A2(\myreg/_1462_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1463_ ) );
AND2_X1 \myreg/_3936_ ( .A1(\myreg/_1457_ ), .A2(\myreg/_1463_ ), .ZN(\myreg/_1464_ ) );
MUX2_X1 \myreg/_3937_ ( .A(\myreg/_0334_ ), .B(\myreg/_0366_ ), .S(fanout_net_35 ), .Z(\myreg/_1465_ ) );
MUX2_X1 \myreg/_3938_ ( .A(\myreg/_0398_ ), .B(\myreg/_0430_ ), .S(fanout_net_35 ), .Z(\myreg/_1466_ ) );
MUX2_X1 \myreg/_3939_ ( .A(\myreg/_1465_ ), .B(\myreg/_1466_ ), .S(fanout_net_42 ), .Z(\myreg/_1467_ ) );
MUX2_X1 \myreg/_3940_ ( .A(\myreg/_0014_ ), .B(\myreg/_0238_ ), .S(fanout_net_35 ), .Z(\myreg/_1468_ ) );
MUX2_X1 \myreg/_3941_ ( .A(\myreg/_0270_ ), .B(\myreg/_0302_ ), .S(fanout_net_35 ), .Z(\myreg/_1469_ ) );
MUX2_X1 \myreg/_3942_ ( .A(\myreg/_1468_ ), .B(\myreg/_1469_ ), .S(fanout_net_42 ), .Z(\myreg/_1470_ ) );
MUX2_X1 \myreg/_3943_ ( .A(\myreg/_1467_ ), .B(\myreg/_1470_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1471_ ) );
MUX2_X1 \myreg/_3944_ ( .A(\myreg/_1464_ ), .B(\myreg/_1471_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2362_ ) );
MUX2_X1 \myreg/_3945_ ( .A(\myreg/_0111_ ), .B(\myreg/_0143_ ), .S(fanout_net_35 ), .Z(\myreg/_1472_ ) );
MUX2_X1 \myreg/_3946_ ( .A(\myreg/_0175_ ), .B(\myreg/_0207_ ), .S(fanout_net_35 ), .Z(\myreg/_1473_ ) );
MUX2_X1 \myreg/_3947_ ( .A(\myreg/_1472_ ), .B(\myreg/_1473_ ), .S(fanout_net_42 ), .Z(\myreg/_1474_ ) );
MUX2_X1 \myreg/_3948_ ( .A(\myreg/_0463_ ), .B(\myreg/_0495_ ), .S(fanout_net_35 ), .Z(\myreg/_1475_ ) );
MUX2_X1 \myreg/_3949_ ( .A(\myreg/_0047_ ), .B(\myreg/_0079_ ), .S(fanout_net_35 ), .Z(\myreg/_1476_ ) );
MUX2_X1 \myreg/_3950_ ( .A(\myreg/_1475_ ), .B(\myreg/_1476_ ), .S(fanout_net_42 ), .Z(\myreg/_1477_ ) );
MUX2_X1 \myreg/_3951_ ( .A(\myreg/_1474_ ), .B(\myreg/_1477_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1478_ ) );
MUX2_X1 \myreg/_3952_ ( .A(\myreg/_0015_ ), .B(\myreg/_0271_ ), .S(fanout_net_42 ), .Z(\myreg/_1479_ ) );
MUX2_X1 \myreg/_3953_ ( .A(\myreg/_0239_ ), .B(\myreg/_0303_ ), .S(fanout_net_42 ), .Z(\myreg/_1480_ ) );
MUX2_X1 \myreg/_3954_ ( .A(\myreg/_1479_ ), .B(\myreg/_1480_ ), .S(fanout_net_35 ), .Z(\myreg/_1481_ ) );
MUX2_X1 \myreg/_3955_ ( .A(\myreg/_0335_ ), .B(\myreg/_0399_ ), .S(fanout_net_42 ), .Z(\myreg/_1482_ ) );
MUX2_X1 \myreg/_3956_ ( .A(\myreg/_0367_ ), .B(\myreg/_0431_ ), .S(fanout_net_42 ), .Z(\myreg/_1483_ ) );
MUX2_X1 \myreg/_3957_ ( .A(\myreg/_1482_ ), .B(\myreg/_1483_ ), .S(fanout_net_35 ), .Z(\myreg/_1484_ ) );
MUX2_X1 \myreg/_3958_ ( .A(\myreg/_1481_ ), .B(\myreg/_1484_ ), .S(fanout_net_44 ), .Z(\myreg/_1485_ ) );
MUX2_X1 \myreg/_3959_ ( .A(\myreg/_1478_ ), .B(\myreg/_1485_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2363_ ) );
NOR2_X1 \myreg/_3960_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0144_ ), .ZN(\myreg/_1486_ ) );
NOR2_X1 \myreg/_3961_ ( .A1(fanout_net_35 ), .A2(\myreg/_0112_ ), .ZN(\myreg/_1487_ ) );
OR3_X1 \myreg/_3962_ ( .A1(\myreg/_1486_ ), .A2(fanout_net_42 ), .A3(\myreg/_1487_ ), .ZN(\myreg/_1488_ ) );
OR2_X1 \myreg/_3963_ ( .A1(\myreg/_1025_ ), .A2(\myreg/_0208_ ), .ZN(\myreg/_1489_ ) );
OAI211_X2 \myreg/_3964_ ( .A(\myreg/_1489_ ), .B(fanout_net_42 ), .C1(fanout_net_36 ), .C2(\myreg/_0176_ ), .ZN(\myreg/_1490_ ) );
AOI21_X1 \myreg/_3965_ ( .A(\myreg/_1039_ ), .B1(\myreg/_1488_ ), .B2(\myreg/_1490_ ), .ZN(\myreg/_1491_ ) );
NOR2_X1 \myreg/_3966_ ( .A1(\myreg/_1025_ ), .A2(\myreg/_0496_ ), .ZN(\myreg/_1492_ ) );
NOR2_X1 \myreg/_3967_ ( .A1(fanout_net_36 ), .A2(\myreg/_0464_ ), .ZN(\myreg/_1493_ ) );
OR3_X1 \myreg/_3968_ ( .A1(\myreg/_1492_ ), .A2(fanout_net_42 ), .A3(\myreg/_1493_ ), .ZN(\myreg/_1494_ ) );
OR2_X1 \myreg/_3969_ ( .A1(fanout_net_36 ), .A2(\myreg/_0048_ ), .ZN(\myreg/_1495_ ) );
OAI211_X2 \myreg/_3970_ ( .A(\myreg/_1495_ ), .B(fanout_net_42 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0080_ ), .ZN(\myreg/_1496_ ) );
AOI21_X1 \myreg/_3971_ ( .A(fanout_net_44 ), .B1(\myreg/_1494_ ), .B2(\myreg/_1496_ ), .ZN(\myreg/_1497_ ) );
OR2_X1 \myreg/_3972_ ( .A1(\myreg/_1491_ ), .A2(\myreg/_1497_ ), .ZN(\myreg/_1498_ ) );
MUX2_X1 \myreg/_3973_ ( .A(\myreg/_0336_ ), .B(\myreg/_0368_ ), .S(fanout_net_36 ), .Z(\myreg/_1499_ ) );
MUX2_X1 \myreg/_3974_ ( .A(\myreg/_0400_ ), .B(\myreg/_0432_ ), .S(fanout_net_36 ), .Z(\myreg/_1500_ ) );
MUX2_X1 \myreg/_3975_ ( .A(\myreg/_1499_ ), .B(\myreg/_1500_ ), .S(fanout_net_42 ), .Z(\myreg/_1501_ ) );
MUX2_X1 \myreg/_3976_ ( .A(\myreg/_0016_ ), .B(\myreg/_0240_ ), .S(fanout_net_36 ), .Z(\myreg/_1502_ ) );
MUX2_X1 \myreg/_3977_ ( .A(\myreg/_0272_ ), .B(\myreg/_0304_ ), .S(fanout_net_36 ), .Z(\myreg/_1503_ ) );
MUX2_X1 \myreg/_3978_ ( .A(\myreg/_1502_ ), .B(\myreg/_1503_ ), .S(fanout_net_42 ), .Z(\myreg/_1504_ ) );
MUX2_X1 \myreg/_3979_ ( .A(\myreg/_1501_ ), .B(\myreg/_1504_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1505_ ) );
MUX2_X1 \myreg/_3980_ ( .A(\myreg/_1498_ ), .B(\myreg/_1505_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2364_ ) );
NOR2_X1 \myreg/_3981_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0145_ ), .ZN(\myreg/_1506_ ) );
NOR2_X1 \myreg/_3982_ ( .A1(fanout_net_36 ), .A2(\myreg/_0113_ ), .ZN(\myreg/_1507_ ) );
OR3_X1 \myreg/_3983_ ( .A1(\myreg/_1506_ ), .A2(fanout_net_43 ), .A3(\myreg/_1507_ ), .ZN(\myreg/_1508_ ) );
OR2_X1 \myreg/_3984_ ( .A1(\myreg/_1025_ ), .A2(\myreg/_0209_ ), .ZN(\myreg/_1509_ ) );
OAI211_X2 \myreg/_3985_ ( .A(\myreg/_1509_ ), .B(fanout_net_43 ), .C1(fanout_net_36 ), .C2(\myreg/_0177_ ), .ZN(\myreg/_1510_ ) );
AOI21_X1 \myreg/_3986_ ( .A(\myreg/_1039_ ), .B1(\myreg/_1508_ ), .B2(\myreg/_1510_ ), .ZN(\myreg/_1511_ ) );
NOR2_X1 \myreg/_3987_ ( .A1(\myreg/_1025_ ), .A2(\myreg/_0497_ ), .ZN(\myreg/_1512_ ) );
NOR2_X1 \myreg/_3988_ ( .A1(fanout_net_36 ), .A2(\myreg/_0465_ ), .ZN(\myreg/_1513_ ) );
OR3_X1 \myreg/_3989_ ( .A1(\myreg/_1512_ ), .A2(fanout_net_43 ), .A3(\myreg/_1513_ ), .ZN(\myreg/_1514_ ) );
OR2_X1 \myreg/_3990_ ( .A1(fanout_net_36 ), .A2(\myreg/_0049_ ), .ZN(\myreg/_1515_ ) );
OAI211_X2 \myreg/_3991_ ( .A(\myreg/_1515_ ), .B(fanout_net_43 ), .C1(\myreg/_1026_ ), .C2(\myreg/_0081_ ), .ZN(\myreg/_1516_ ) );
AOI21_X1 \myreg/_3992_ ( .A(fanout_net_44 ), .B1(\myreg/_1514_ ), .B2(\myreg/_1516_ ), .ZN(\myreg/_1517_ ) );
OR2_X1 \myreg/_3993_ ( .A1(\myreg/_1511_ ), .A2(\myreg/_1517_ ), .ZN(\myreg/_1518_ ) );
MUX2_X1 \myreg/_3994_ ( .A(\myreg/_0337_ ), .B(\myreg/_0369_ ), .S(fanout_net_36 ), .Z(\myreg/_1519_ ) );
MUX2_X1 \myreg/_3995_ ( .A(\myreg/_0401_ ), .B(\myreg/_0433_ ), .S(fanout_net_36 ), .Z(\myreg/_1520_ ) );
MUX2_X1 \myreg/_3996_ ( .A(\myreg/_1519_ ), .B(\myreg/_1520_ ), .S(fanout_net_43 ), .Z(\myreg/_1521_ ) );
MUX2_X1 \myreg/_3997_ ( .A(\myreg/_0017_ ), .B(\myreg/_0241_ ), .S(fanout_net_36 ), .Z(\myreg/_1522_ ) );
MUX2_X1 \myreg/_3998_ ( .A(\myreg/_0273_ ), .B(\myreg/_0305_ ), .S(fanout_net_36 ), .Z(\myreg/_1523_ ) );
MUX2_X1 \myreg/_3999_ ( .A(\myreg/_1522_ ), .B(\myreg/_1523_ ), .S(fanout_net_43 ), .Z(\myreg/_1524_ ) );
MUX2_X1 \myreg/_4000_ ( .A(\myreg/_1521_ ), .B(\myreg/_1524_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1525_ ) );
MUX2_X1 \myreg/_4001_ ( .A(\myreg/_1518_ ), .B(\myreg/_1525_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2365_ ) );
OR2_X1 \myreg/_4002_ ( .A1(fanout_net_36 ), .A2(\myreg/_0178_ ), .ZN(\myreg/_1526_ ) );
OAI211_X2 \myreg/_4003_ ( .A(\myreg/_1526_ ), .B(fanout_net_43 ), .C1(\myreg/_1027_ ), .C2(\myreg/_0210_ ), .ZN(\myreg/_1527_ ) );
INV_X1 \myreg/_4004_ ( .A(\myreg/_0146_ ), .ZN(\myreg/_1528_ ) );
AOI21_X1 \myreg/_4005_ ( .A(fanout_net_43 ), .B1(\myreg/_1528_ ), .B2(fanout_net_36 ), .ZN(\myreg/_1529_ ) );
OAI21_X1 \myreg/_4006_ ( .A(\myreg/_1529_ ), .B1(fanout_net_36 ), .B2(\myreg/_0114_ ), .ZN(\myreg/_1530_ ) );
NAND3_X1 \myreg/_4007_ ( .A1(\myreg/_1527_ ), .A2(\myreg/_1530_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1531_ ) );
OR2_X1 \myreg/_4008_ ( .A1(fanout_net_36 ), .A2(\myreg/_0050_ ), .ZN(\myreg/_1532_ ) );
OAI211_X2 \myreg/_4009_ ( .A(\myreg/_1532_ ), .B(fanout_net_43 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0082_ ), .ZN(\myreg/_1533_ ) );
INV_X1 \myreg/_4010_ ( .A(\myreg/_0498_ ), .ZN(\myreg/_1534_ ) );
AOI21_X1 \myreg/_4011_ ( .A(fanout_net_43 ), .B1(\myreg/_1534_ ), .B2(fanout_net_36 ), .ZN(\myreg/_1535_ ) );
OAI21_X1 \myreg/_4012_ ( .A(\myreg/_1535_ ), .B1(fanout_net_36 ), .B2(\myreg/_0466_ ), .ZN(\myreg/_1536_ ) );
NAND3_X1 \myreg/_4013_ ( .A1(\myreg/_1533_ ), .A2(\myreg/_1536_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1537_ ) );
AND2_X1 \myreg/_4014_ ( .A1(\myreg/_1531_ ), .A2(\myreg/_1537_ ), .ZN(\myreg/_1538_ ) );
MUX2_X1 \myreg/_4015_ ( .A(\myreg/_0338_ ), .B(\myreg/_0370_ ), .S(fanout_net_36 ), .Z(\myreg/_1539_ ) );
MUX2_X1 \myreg/_4016_ ( .A(\myreg/_0402_ ), .B(\myreg/_0434_ ), .S(fanout_net_36 ), .Z(\myreg/_1540_ ) );
MUX2_X1 \myreg/_4017_ ( .A(\myreg/_1539_ ), .B(\myreg/_1540_ ), .S(fanout_net_43 ), .Z(\myreg/_1541_ ) );
MUX2_X1 \myreg/_4018_ ( .A(\myreg/_0018_ ), .B(\myreg/_0242_ ), .S(fanout_net_36 ), .Z(\myreg/_1542_ ) );
MUX2_X1 \myreg/_4019_ ( .A(\myreg/_0274_ ), .B(\myreg/_0306_ ), .S(fanout_net_36 ), .Z(\myreg/_1543_ ) );
MUX2_X1 \myreg/_4020_ ( .A(\myreg/_1542_ ), .B(\myreg/_1543_ ), .S(fanout_net_43 ), .Z(\myreg/_1544_ ) );
MUX2_X1 \myreg/_4021_ ( .A(\myreg/_1541_ ), .B(\myreg/_1544_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1545_ ) );
MUX2_X1 \myreg/_4022_ ( .A(\myreg/_1538_ ), .B(\myreg/_1545_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2366_ ) );
OR2_X1 \myreg/_4023_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0083_ ), .ZN(\myreg/_1546_ ) );
OAI211_X2 \myreg/_4024_ ( .A(\myreg/_1546_ ), .B(fanout_net_43 ), .C1(fanout_net_36 ), .C2(\myreg/_0051_ ), .ZN(\myreg/_1547_ ) );
INV_X1 \myreg/_4025_ ( .A(\myreg/_0499_ ), .ZN(\myreg/_1548_ ) );
AOI21_X1 \myreg/_4026_ ( .A(fanout_net_43 ), .B1(\myreg/_1548_ ), .B2(fanout_net_36 ), .ZN(\myreg/_1549_ ) );
OAI21_X1 \myreg/_4027_ ( .A(\myreg/_1549_ ), .B1(fanout_net_36 ), .B2(\myreg/_0467_ ), .ZN(\myreg/_1550_ ) );
NAND3_X1 \myreg/_4028_ ( .A1(\myreg/_1547_ ), .A2(\myreg/_1040_ ), .A3(\myreg/_1550_ ), .ZN(\myreg/_1551_ ) );
OR2_X1 \myreg/_4029_ ( .A1(fanout_net_36 ), .A2(\myreg/_0179_ ), .ZN(\myreg/_1552_ ) );
OAI211_X2 \myreg/_4030_ ( .A(\myreg/_1552_ ), .B(fanout_net_43 ), .C1(\myreg/_1227_ ), .C2(\myreg/_0211_ ), .ZN(\myreg/_1553_ ) );
INV_X1 \myreg/_4031_ ( .A(\myreg/_0147_ ), .ZN(\myreg/_1554_ ) );
AOI21_X1 \myreg/_4032_ ( .A(fanout_net_43 ), .B1(\myreg/_1554_ ), .B2(fanout_net_36 ), .ZN(\myreg/_1555_ ) );
OAI21_X1 \myreg/_4033_ ( .A(\myreg/_1555_ ), .B1(fanout_net_37 ), .B2(\myreg/_0115_ ), .ZN(\myreg/_1556_ ) );
NAND3_X1 \myreg/_4034_ ( .A1(\myreg/_1553_ ), .A2(\myreg/_1556_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1557_ ) );
AND2_X1 \myreg/_4035_ ( .A1(\myreg/_1551_ ), .A2(\myreg/_1557_ ), .ZN(\myreg/_1558_ ) );
MUX2_X1 \myreg/_4036_ ( .A(\myreg/_0339_ ), .B(\myreg/_0371_ ), .S(fanout_net_37 ), .Z(\myreg/_1559_ ) );
MUX2_X1 \myreg/_4037_ ( .A(\myreg/_0403_ ), .B(\myreg/_0435_ ), .S(fanout_net_37 ), .Z(\myreg/_1560_ ) );
MUX2_X1 \myreg/_4038_ ( .A(\myreg/_1559_ ), .B(\myreg/_1560_ ), .S(fanout_net_43 ), .Z(\myreg/_1561_ ) );
MUX2_X1 \myreg/_4039_ ( .A(\myreg/_0019_ ), .B(\myreg/_0243_ ), .S(fanout_net_37 ), .Z(\myreg/_1562_ ) );
MUX2_X1 \myreg/_4040_ ( .A(\myreg/_0275_ ), .B(\myreg/_0307_ ), .S(fanout_net_37 ), .Z(\myreg/_1563_ ) );
MUX2_X1 \myreg/_4041_ ( .A(\myreg/_1562_ ), .B(\myreg/_1563_ ), .S(fanout_net_43 ), .Z(\myreg/_1564_ ) );
MUX2_X1 \myreg/_4042_ ( .A(\myreg/_1561_ ), .B(\myreg/_1564_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1565_ ) );
MUX2_X1 \myreg/_4043_ ( .A(\myreg/_1558_ ), .B(\myreg/_1565_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2367_ ) );
NOR2_X1 \myreg/_4044_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0148_ ), .ZN(\myreg/_1566_ ) );
NOR2_X1 \myreg/_4045_ ( .A1(fanout_net_37 ), .A2(\myreg/_0116_ ), .ZN(\myreg/_1567_ ) );
OR3_X1 \myreg/_4046_ ( .A1(\myreg/_1566_ ), .A2(fanout_net_43 ), .A3(\myreg/_1567_ ), .ZN(\myreg/_1568_ ) );
OR2_X1 \myreg/_4047_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0212_ ), .ZN(\myreg/_1569_ ) );
OAI211_X2 \myreg/_4048_ ( .A(\myreg/_1569_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg/_0180_ ), .ZN(\myreg/_1570_ ) );
NAND3_X1 \myreg/_4049_ ( .A1(\myreg/_1568_ ), .A2(\myreg/_1570_ ), .A3(fanout_net_44 ), .ZN(\myreg/_1571_ ) );
NOR2_X1 \myreg/_4050_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0500_ ), .ZN(\myreg/_1572_ ) );
NOR2_X1 \myreg/_4051_ ( .A1(fanout_net_37 ), .A2(\myreg/_0468_ ), .ZN(\myreg/_1573_ ) );
OR3_X1 \myreg/_4052_ ( .A1(\myreg/_1572_ ), .A2(fanout_net_43 ), .A3(\myreg/_1573_ ), .ZN(\myreg/_1574_ ) );
OR2_X1 \myreg/_4053_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0084_ ), .ZN(\myreg/_1575_ ) );
OAI211_X2 \myreg/_4054_ ( .A(\myreg/_1575_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg/_0052_ ), .ZN(\myreg/_1576_ ) );
NAND3_X1 \myreg/_4055_ ( .A1(\myreg/_1574_ ), .A2(\myreg/_1576_ ), .A3(\myreg/_1049_ ), .ZN(\myreg/_1577_ ) );
AND2_X1 \myreg/_4056_ ( .A1(\myreg/_1571_ ), .A2(\myreg/_1577_ ), .ZN(\myreg/_1578_ ) );
MUX2_X1 \myreg/_4057_ ( .A(\myreg/_0340_ ), .B(\myreg/_0372_ ), .S(fanout_net_37 ), .Z(\myreg/_1579_ ) );
MUX2_X1 \myreg/_4058_ ( .A(\myreg/_0404_ ), .B(\myreg/_0436_ ), .S(fanout_net_37 ), .Z(\myreg/_1580_ ) );
MUX2_X1 \myreg/_4059_ ( .A(\myreg/_1579_ ), .B(\myreg/_1580_ ), .S(fanout_net_43 ), .Z(\myreg/_1581_ ) );
MUX2_X1 \myreg/_4060_ ( .A(\myreg/_0020_ ), .B(\myreg/_0244_ ), .S(fanout_net_37 ), .Z(\myreg/_1582_ ) );
MUX2_X1 \myreg/_4061_ ( .A(\myreg/_0276_ ), .B(\myreg/_0308_ ), .S(fanout_net_37 ), .Z(\myreg/_1583_ ) );
MUX2_X1 \myreg/_4062_ ( .A(\myreg/_1582_ ), .B(\myreg/_1583_ ), .S(fanout_net_43 ), .Z(\myreg/_1584_ ) );
MUX2_X1 \myreg/_4063_ ( .A(\myreg/_1581_ ), .B(\myreg/_1584_ ), .S(\myreg/_1389_ ), .Z(\myreg/_1585_ ) );
MUX2_X1 \myreg/_4064_ ( .A(\myreg/_1578_ ), .B(\myreg/_1585_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2368_ ) );
NOR2_X1 \myreg/_4065_ ( .A1(\myreg/_1026_ ), .A2(\myreg/_0501_ ), .ZN(\myreg/_1586_ ) );
NOR2_X1 \myreg/_4066_ ( .A1(fanout_net_37 ), .A2(\myreg/_0469_ ), .ZN(\myreg/_1587_ ) );
OR3_X1 \myreg/_4067_ ( .A1(\myreg/_1586_ ), .A2(fanout_net_43 ), .A3(\myreg/_1587_ ), .ZN(\myreg/_1588_ ) );
OR2_X1 \myreg/_4068_ ( .A1(\myreg/_1199_ ), .A2(\myreg/_0085_ ), .ZN(\myreg/_1589_ ) );
OAI211_X2 \myreg/_4069_ ( .A(\myreg/_1589_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg/_0053_ ), .ZN(\myreg/_1590_ ) );
NAND3_X1 \myreg/_4070_ ( .A1(\myreg/_1588_ ), .A2(\myreg/_1590_ ), .A3(\myreg/_1040_ ), .ZN(\myreg/_1591_ ) );
NOR2_X1 \myreg/_4071_ ( .A1(\myreg/_1074_ ), .A2(\myreg/_0149_ ), .ZN(\myreg/_1592_ ) );
NOR2_X1 \myreg/_4072_ ( .A1(fanout_net_37 ), .A2(\myreg/_0117_ ), .ZN(\myreg/_1593_ ) );
OR3_X1 \myreg/_4073_ ( .A1(\myreg/_1592_ ), .A2(fanout_net_43 ), .A3(\myreg/_1593_ ), .ZN(\myreg/_1594_ ) );
OR2_X1 \myreg/_4074_ ( .A1(fanout_net_37 ), .A2(\myreg/_0181_ ), .ZN(\myreg/_1595_ ) );
OAI211_X2 \myreg/_4075_ ( .A(\myreg/_1595_ ), .B(fanout_net_43 ), .C1(\myreg/_1054_ ), .C2(\myreg/_0213_ ), .ZN(\myreg/_1596_ ) );
NAND3_X1 \myreg/_4076_ ( .A1(\myreg/_1594_ ), .A2(\myreg/_2342_ ), .A3(\myreg/_1596_ ), .ZN(\myreg/_1597_ ) );
AND2_X1 \myreg/_4077_ ( .A1(\myreg/_1591_ ), .A2(\myreg/_1597_ ), .ZN(\myreg/_1598_ ) );
MUX2_X1 \myreg/_4078_ ( .A(\myreg/_0341_ ), .B(\myreg/_0373_ ), .S(fanout_net_37 ), .Z(\myreg/_1599_ ) );
MUX2_X1 \myreg/_4079_ ( .A(\myreg/_0405_ ), .B(\myreg/_0437_ ), .S(fanout_net_37 ), .Z(\myreg/_1600_ ) );
MUX2_X1 \myreg/_4080_ ( .A(\myreg/_1599_ ), .B(\myreg/_1600_ ), .S(fanout_net_43 ), .Z(\myreg/_1601_ ) );
MUX2_X1 \myreg/_4081_ ( .A(\myreg/_0021_ ), .B(\myreg/_0245_ ), .S(fanout_net_37 ), .Z(\myreg/_1602_ ) );
MUX2_X1 \myreg/_4082_ ( .A(\myreg/_0277_ ), .B(\myreg/_0309_ ), .S(fanout_net_37 ), .Z(\myreg/_1603_ ) );
MUX2_X1 \myreg/_4083_ ( .A(\myreg/_1602_ ), .B(\myreg/_1603_ ), .S(fanout_net_43 ), .Z(\myreg/_1604_ ) );
MUX2_X1 \myreg/_4084_ ( .A(\myreg/_1601_ ), .B(\myreg/_1604_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1605_ ) );
MUX2_X1 \myreg/_4085_ ( .A(\myreg/_1598_ ), .B(\myreg/_1605_ ), .S(\myreg/_1431_ ), .Z(\myreg/_2369_ ) );
MUX2_X1 \myreg/_4086_ ( .A(\myreg/_0119_ ), .B(\myreg/_0151_ ), .S(fanout_net_37 ), .Z(\myreg/_1606_ ) );
MUX2_X1 \myreg/_4087_ ( .A(\myreg/_0183_ ), .B(\myreg/_0215_ ), .S(fanout_net_37 ), .Z(\myreg/_1607_ ) );
MUX2_X1 \myreg/_4088_ ( .A(\myreg/_1606_ ), .B(\myreg/_1607_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1608_ ) );
MUX2_X1 \myreg/_4089_ ( .A(\myreg/_0471_ ), .B(\myreg/_0503_ ), .S(fanout_net_37 ), .Z(\myreg/_1609_ ) );
MUX2_X1 \myreg/_4090_ ( .A(\myreg/_0055_ ), .B(\myreg/_0087_ ), .S(fanout_net_37 ), .Z(\myreg/_1610_ ) );
MUX2_X1 \myreg/_4091_ ( .A(\myreg/_1609_ ), .B(\myreg/_1610_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1611_ ) );
MUX2_X1 \myreg/_4092_ ( .A(\myreg/_1608_ ), .B(\myreg/_1611_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1612_ ) );
MUX2_X1 \myreg/_4093_ ( .A(\myreg/_0023_ ), .B(\myreg/_0279_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1613_ ) );
MUX2_X1 \myreg/_4094_ ( .A(\myreg/_0247_ ), .B(\myreg/_0311_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1614_ ) );
MUX2_X1 \myreg/_4095_ ( .A(\myreg/_1613_ ), .B(\myreg/_1614_ ), .S(fanout_net_37 ), .Z(\myreg/_1615_ ) );
MUX2_X1 \myreg/_4096_ ( .A(\myreg/_0343_ ), .B(\myreg/_0407_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1616_ ) );
MUX2_X1 \myreg/_4097_ ( .A(\myreg/_0375_ ), .B(\myreg/_0439_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1617_ ) );
MUX2_X1 \myreg/_4098_ ( .A(\myreg/_1616_ ), .B(\myreg/_1617_ ), .S(fanout_net_37 ), .Z(\myreg/_1618_ ) );
MUX2_X1 \myreg/_4099_ ( .A(\myreg/_1615_ ), .B(\myreg/_1618_ ), .S(\myreg/_2342_ ), .Z(\myreg/_1619_ ) );
MUX2_X1 \myreg/_4100_ ( .A(\myreg/_1612_ ), .B(\myreg/_1619_ ), .S(\myreg/_1051_ ), .Z(\myreg/_2371_ ) );
MUX2_X1 \myreg/_4101_ ( .A(\myreg/_0120_ ), .B(\myreg/_0152_ ), .S(fanout_net_37 ), .Z(\myreg/_1620_ ) );
MUX2_X1 \myreg/_4102_ ( .A(\myreg/_0184_ ), .B(\myreg/_0216_ ), .S(fanout_net_37 ), .Z(\myreg/_1621_ ) );
MUX2_X1 \myreg/_4103_ ( .A(\myreg/_1620_ ), .B(\myreg/_1621_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1622_ ) );
MUX2_X1 \myreg/_4104_ ( .A(\myreg/_0472_ ), .B(\myreg/_0504_ ), .S(fanout_net_37 ), .Z(\myreg/_1623_ ) );
MUX2_X1 \myreg/_4105_ ( .A(\myreg/_0056_ ), .B(\myreg/_0088_ ), .S(\myreg/_2340_ ), .Z(\myreg/_1624_ ) );
MUX2_X1 \myreg/_4106_ ( .A(\myreg/_1623_ ), .B(\myreg/_1624_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1625_ ) );
MUX2_X1 \myreg/_4107_ ( .A(\myreg/_1622_ ), .B(\myreg/_1625_ ), .S(\myreg/_1142_ ), .Z(\myreg/_1626_ ) );
MUX2_X1 \myreg/_4108_ ( .A(\myreg/_0024_ ), .B(\myreg/_0280_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1627_ ) );
MUX2_X1 \myreg/_4109_ ( .A(\myreg/_0248_ ), .B(\myreg/_0312_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1628_ ) );
MUX2_X1 \myreg/_4110_ ( .A(\myreg/_1627_ ), .B(\myreg/_1628_ ), .S(\myreg/_2340_ ), .Z(\myreg/_1629_ ) );
MUX2_X1 \myreg/_4111_ ( .A(\myreg/_0344_ ), .B(\myreg/_0408_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1630_ ) );
MUX2_X1 \myreg/_4112_ ( .A(\myreg/_0376_ ), .B(\myreg/_0440_ ), .S(\myreg/_2341_ ), .Z(\myreg/_1631_ ) );
MUX2_X1 \myreg/_4113_ ( .A(\myreg/_1630_ ), .B(\myreg/_1631_ ), .S(\myreg/_2340_ ), .Z(\myreg/_1632_ ) );
MUX2_X1 \myreg/_4114_ ( .A(\myreg/_1629_ ), .B(\myreg/_1632_ ), .S(\myreg/_2342_ ), .Z(\myreg/_1633_ ) );
MUX2_X1 \myreg/_4115_ ( .A(\myreg/_1626_ ), .B(\myreg/_1633_ ), .S(\myreg/_1051_ ), .Z(\myreg/_2372_ ) );
INV_X1 \myreg/_4116_ ( .A(fanout_net_45 ), .ZN(\myreg/_1634_ ) );
BUF_X2 \myreg/_4117_ ( .A(\myreg/_1634_ ), .Z(\myreg/_1635_ ) );
OR2_X1 \myreg/_4118_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0064_ ), .ZN(\myreg/_1636_ ) );
OAI211_X2 \myreg/_4119_ ( .A(\myreg/_1636_ ), .B(fanout_net_54 ), .C1(\myreg/_0032_ ), .C2(fanout_net_45 ), .ZN(\myreg/_1637_ ) );
AOI21_X1 \myreg/_4120_ ( .A(fanout_net_54 ), .B1(\myreg/_1035_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1638_ ) );
OAI21_X1 \myreg/_4121_ ( .A(\myreg/_1638_ ), .B1(\myreg/_0448_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1639_ ) );
AOI21_X1 \myreg/_4122_ ( .A(fanout_net_60 ), .B1(\myreg/_1637_ ), .B2(\myreg/_1639_ ), .ZN(\myreg/_1640_ ) );
INV_X1 \myreg/_4123_ ( .A(fanout_net_60 ), .ZN(\myreg/_1641_ ) );
BUF_X4 \myreg/_4124_ ( .A(\myreg/_1641_ ), .Z(\myreg/_1642_ ) );
OR2_X1 \myreg/_4125_ ( .A1(\myreg/_0160_ ), .A2(fanout_net_45 ), .ZN(\myreg/_1643_ ) );
BUF_X8 \myreg/_4126_ ( .A(\myreg/_1635_ ), .Z(\myreg/_1644_ ) );
OAI211_X2 \myreg/_4127_ ( .A(\myreg/_1643_ ), .B(fanout_net_54 ), .C1(\myreg/_0192_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1645_ ) );
AOI21_X1 \myreg/_4128_ ( .A(fanout_net_54 ), .B1(\myreg/_1029_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1646_ ) );
OAI21_X1 \myreg/_4129_ ( .A(\myreg/_1646_ ), .B1(\myreg/_0096_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1647_ ) );
AOI21_X1 \myreg/_4130_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1645_ ), .B2(\myreg/_1647_ ), .ZN(\myreg/_1648_ ) );
OR2_X1 \myreg/_4131_ ( .A1(\myreg/_1640_ ), .A2(\myreg/_1648_ ), .ZN(\myreg/_1649_ ) );
MUX2_X1 \myreg/_4132_ ( .A(\myreg/_0320_ ), .B(\myreg/_0352_ ), .S(fanout_net_45 ), .Z(\myreg/_1650_ ) );
MUX2_X1 \myreg/_4133_ ( .A(\myreg/_0384_ ), .B(\myreg/_0416_ ), .S(fanout_net_45 ), .Z(\myreg/_1651_ ) );
MUX2_X1 \myreg/_4134_ ( .A(\myreg/_1650_ ), .B(\myreg/_1651_ ), .S(fanout_net_54 ), .Z(\myreg/_1652_ ) );
MUX2_X1 \myreg/_4135_ ( .A(\myreg/_0000_ ), .B(\myreg/_0224_ ), .S(fanout_net_45 ), .Z(\myreg/_1653_ ) );
MUX2_X1 \myreg/_4136_ ( .A(\myreg/_0256_ ), .B(\myreg/_0288_ ), .S(fanout_net_45 ), .Z(\myreg/_1654_ ) );
MUX2_X1 \myreg/_4137_ ( .A(\myreg/_1653_ ), .B(\myreg/_1654_ ), .S(fanout_net_54 ), .Z(\myreg/_1655_ ) );
BUF_X4 \myreg/_4138_ ( .A(\myreg/_1642_ ), .Z(\myreg/_1656_ ) );
MUX2_X1 \myreg/_4139_ ( .A(\myreg/_1652_ ), .B(\myreg/_1655_ ), .S(\myreg/_1656_ ), .Z(\myreg/_1657_ ) );
INV_X1 \myreg/_4140_ ( .A(\myreg/_2347_ ), .ZN(\myreg/_1658_ ) );
BUF_X4 \myreg/_4141_ ( .A(\myreg/_1658_ ), .Z(\myreg/_1659_ ) );
MUX2_X1 \myreg/_4142_ ( .A(\myreg/_1649_ ), .B(\myreg/_1657_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2380_ ) );
BUF_X4 \myreg/_4143_ ( .A(\myreg/_1641_ ), .Z(\myreg/_1660_ ) );
OR2_X1 \myreg/_4144_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0203_ ), .ZN(\myreg/_1661_ ) );
OAI211_X2 \myreg/_4145_ ( .A(\myreg/_1661_ ), .B(fanout_net_54 ), .C1(\myreg/_0171_ ), .C2(fanout_net_45 ), .ZN(\myreg/_1662_ ) );
AOI21_X1 \myreg/_4146_ ( .A(fanout_net_54 ), .B1(\myreg/_1062_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1663_ ) );
OAI21_X1 \myreg/_4147_ ( .A(\myreg/_1663_ ), .B1(\myreg/_0107_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1664_ ) );
AOI21_X1 \myreg/_4148_ ( .A(\myreg/_1660_ ), .B1(\myreg/_1662_ ), .B2(\myreg/_1664_ ), .ZN(\myreg/_1665_ ) );
OR2_X1 \myreg/_4149_ ( .A1(\myreg/_0043_ ), .A2(fanout_net_45 ), .ZN(\myreg/_1666_ ) );
OAI211_X2 \myreg/_4150_ ( .A(\myreg/_1666_ ), .B(fanout_net_54 ), .C1(\myreg/_0075_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1667_ ) );
AOI21_X1 \myreg/_4151_ ( .A(fanout_net_54 ), .B1(\myreg/_1056_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1668_ ) );
OAI21_X1 \myreg/_4152_ ( .A(\myreg/_1668_ ), .B1(\myreg/_0459_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1669_ ) );
AOI21_X1 \myreg/_4153_ ( .A(fanout_net_60 ), .B1(\myreg/_1667_ ), .B2(\myreg/_1669_ ), .ZN(\myreg/_1670_ ) );
OR2_X1 \myreg/_4154_ ( .A1(\myreg/_1665_ ), .A2(\myreg/_1670_ ), .ZN(\myreg/_1671_ ) );
MUX2_X1 \myreg/_4155_ ( .A(\myreg/_0331_ ), .B(\myreg/_0363_ ), .S(fanout_net_45 ), .Z(\myreg/_1672_ ) );
MUX2_X1 \myreg/_4156_ ( .A(\myreg/_0395_ ), .B(\myreg/_0427_ ), .S(fanout_net_45 ), .Z(\myreg/_1673_ ) );
MUX2_X1 \myreg/_4157_ ( .A(\myreg/_1672_ ), .B(\myreg/_1673_ ), .S(fanout_net_54 ), .Z(\myreg/_1674_ ) );
MUX2_X1 \myreg/_4158_ ( .A(\myreg/_0011_ ), .B(\myreg/_0235_ ), .S(fanout_net_45 ), .Z(\myreg/_1675_ ) );
MUX2_X1 \myreg/_4159_ ( .A(\myreg/_0267_ ), .B(\myreg/_0299_ ), .S(fanout_net_45 ), .Z(\myreg/_1676_ ) );
MUX2_X1 \myreg/_4160_ ( .A(\myreg/_1675_ ), .B(\myreg/_1676_ ), .S(fanout_net_54 ), .Z(\myreg/_1677_ ) );
MUX2_X1 \myreg/_4161_ ( .A(\myreg/_1674_ ), .B(\myreg/_1677_ ), .S(\myreg/_1656_ ), .Z(\myreg/_1678_ ) );
MUX2_X1 \myreg/_4162_ ( .A(\myreg/_1671_ ), .B(\myreg/_1678_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2391_ ) );
BUF_X4 \myreg/_4163_ ( .A(\myreg/_1634_ ), .Z(\myreg/_1679_ ) );
OR2_X1 \myreg/_4164_ ( .A1(\myreg/_1679_ ), .A2(\myreg/_0214_ ), .ZN(\myreg/_1680_ ) );
OAI211_X2 \myreg/_4165_ ( .A(\myreg/_1680_ ), .B(fanout_net_54 ), .C1(\myreg/_0182_ ), .C2(fanout_net_45 ), .ZN(\myreg/_1681_ ) );
AOI21_X1 \myreg/_4166_ ( .A(fanout_net_54 ), .B1(\myreg/_1083_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1682_ ) );
OAI21_X1 \myreg/_4167_ ( .A(\myreg/_1682_ ), .B1(\myreg/_0118_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1683_ ) );
NAND3_X1 \myreg/_4168_ ( .A1(\myreg/_1681_ ), .A2(fanout_net_60 ), .A3(\myreg/_1683_ ), .ZN(\myreg/_1684_ ) );
OR2_X1 \myreg/_4169_ ( .A1(\myreg/_0054_ ), .A2(fanout_net_45 ), .ZN(\myreg/_1685_ ) );
OAI211_X2 \myreg/_4170_ ( .A(\myreg/_1685_ ), .B(fanout_net_54 ), .C1(\myreg/_0086_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1686_ ) );
AOI21_X1 \myreg/_4171_ ( .A(fanout_net_54 ), .B1(\myreg/_1077_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1687_ ) );
OAI21_X1 \myreg/_4172_ ( .A(\myreg/_1687_ ), .B1(\myreg/_0470_ ), .B2(fanout_net_45 ), .ZN(\myreg/_1688_ ) );
NAND3_X1 \myreg/_4173_ ( .A1(\myreg/_1686_ ), .A2(\myreg/_1688_ ), .A3(\myreg/_1656_ ), .ZN(\myreg/_1689_ ) );
AND2_X1 \myreg/_4174_ ( .A1(\myreg/_1684_ ), .A2(\myreg/_1689_ ), .ZN(\myreg/_1690_ ) );
MUX2_X1 \myreg/_4175_ ( .A(\myreg/_0342_ ), .B(\myreg/_0374_ ), .S(fanout_net_45 ), .Z(\myreg/_1691_ ) );
MUX2_X1 \myreg/_4176_ ( .A(\myreg/_0406_ ), .B(\myreg/_0438_ ), .S(fanout_net_45 ), .Z(\myreg/_1692_ ) );
MUX2_X1 \myreg/_4177_ ( .A(\myreg/_1691_ ), .B(\myreg/_1692_ ), .S(fanout_net_54 ), .Z(\myreg/_1693_ ) );
MUX2_X1 \myreg/_4178_ ( .A(\myreg/_0022_ ), .B(\myreg/_0246_ ), .S(fanout_net_45 ), .Z(\myreg/_1694_ ) );
MUX2_X1 \myreg/_4179_ ( .A(\myreg/_0278_ ), .B(\myreg/_0310_ ), .S(fanout_net_46 ), .Z(\myreg/_1695_ ) );
MUX2_X1 \myreg/_4180_ ( .A(\myreg/_1694_ ), .B(\myreg/_1695_ ), .S(fanout_net_54 ), .Z(\myreg/_1696_ ) );
MUX2_X1 \myreg/_4181_ ( .A(\myreg/_1693_ ), .B(\myreg/_1696_ ), .S(\myreg/_1656_ ), .Z(\myreg/_1697_ ) );
MUX2_X1 \myreg/_4182_ ( .A(\myreg/_1690_ ), .B(\myreg/_1697_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2402_ ) );
OR2_X1 \myreg/_4183_ ( .A1(\myreg/_1679_ ), .A2(\myreg/_0089_ ), .ZN(\myreg/_1698_ ) );
OAI211_X2 \myreg/_4184_ ( .A(\myreg/_1698_ ), .B(fanout_net_54 ), .C1(\myreg/_0057_ ), .C2(fanout_net_46 ), .ZN(\myreg/_1699_ ) );
AOI21_X1 \myreg/_4185_ ( .A(fanout_net_54 ), .B1(\myreg/_1103_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1700_ ) );
OAI21_X1 \myreg/_4186_ ( .A(\myreg/_1700_ ), .B1(\myreg/_0473_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1701_ ) );
NAND3_X1 \myreg/_4187_ ( .A1(\myreg/_1699_ ), .A2(\myreg/_1656_ ), .A3(\myreg/_1701_ ), .ZN(\myreg/_1702_ ) );
OR2_X1 \myreg/_4188_ ( .A1(\myreg/_0185_ ), .A2(fanout_net_46 ), .ZN(\myreg/_1703_ ) );
OAI211_X2 \myreg/_4189_ ( .A(\myreg/_1703_ ), .B(fanout_net_54 ), .C1(\myreg/_0217_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1704_ ) );
AOI21_X1 \myreg/_4190_ ( .A(fanout_net_54 ), .B1(\myreg/_1097_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1705_ ) );
OAI21_X1 \myreg/_4191_ ( .A(\myreg/_1705_ ), .B1(\myreg/_0121_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1706_ ) );
NAND3_X1 \myreg/_4192_ ( .A1(\myreg/_1704_ ), .A2(\myreg/_1706_ ), .A3(fanout_net_60 ), .ZN(\myreg/_1707_ ) );
AND2_X1 \myreg/_4193_ ( .A1(\myreg/_1702_ ), .A2(\myreg/_1707_ ), .ZN(\myreg/_1708_ ) );
MUX2_X1 \myreg/_4194_ ( .A(\myreg/_0345_ ), .B(\myreg/_0377_ ), .S(fanout_net_46 ), .Z(\myreg/_1709_ ) );
MUX2_X1 \myreg/_4195_ ( .A(\myreg/_0409_ ), .B(\myreg/_0441_ ), .S(fanout_net_46 ), .Z(\myreg/_1710_ ) );
MUX2_X1 \myreg/_4196_ ( .A(\myreg/_1709_ ), .B(\myreg/_1710_ ), .S(fanout_net_54 ), .Z(\myreg/_1711_ ) );
MUX2_X1 \myreg/_4197_ ( .A(\myreg/_0025_ ), .B(\myreg/_0249_ ), .S(fanout_net_46 ), .Z(\myreg/_1712_ ) );
MUX2_X1 \myreg/_4198_ ( .A(\myreg/_0281_ ), .B(\myreg/_0313_ ), .S(fanout_net_46 ), .Z(\myreg/_1713_ ) );
MUX2_X1 \myreg/_4199_ ( .A(\myreg/_1712_ ), .B(\myreg/_1713_ ), .S(fanout_net_54 ), .Z(\myreg/_1714_ ) );
BUF_X4 \myreg/_4200_ ( .A(\myreg/_1642_ ), .Z(\myreg/_1715_ ) );
MUX2_X1 \myreg/_4201_ ( .A(\myreg/_1711_ ), .B(\myreg/_1714_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1716_ ) );
MUX2_X1 \myreg/_4202_ ( .A(\myreg/_1708_ ), .B(\myreg/_1716_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2405_ ) );
OR2_X1 \myreg/_4203_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0090_ ), .ZN(\myreg/_1717_ ) );
OAI211_X2 \myreg/_4204_ ( .A(\myreg/_1717_ ), .B(fanout_net_54 ), .C1(\myreg/_0058_ ), .C2(fanout_net_46 ), .ZN(\myreg/_1718_ ) );
AOI21_X1 \myreg/_4205_ ( .A(fanout_net_54 ), .B1(\myreg/_1124_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1719_ ) );
OAI21_X1 \myreg/_4206_ ( .A(\myreg/_1719_ ), .B1(\myreg/_0474_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1720_ ) );
AOI21_X1 \myreg/_4207_ ( .A(fanout_net_60 ), .B1(\myreg/_1718_ ), .B2(\myreg/_1720_ ), .ZN(\myreg/_1721_ ) );
OR2_X1 \myreg/_4208_ ( .A1(\myreg/_1634_ ), .A2(\myreg/_0218_ ), .ZN(\myreg/_1722_ ) );
OAI211_X2 \myreg/_4209_ ( .A(\myreg/_1722_ ), .B(fanout_net_54 ), .C1(\myreg/_0186_ ), .C2(fanout_net_46 ), .ZN(\myreg/_1723_ ) );
AOI21_X1 \myreg/_4210_ ( .A(fanout_net_54 ), .B1(\myreg/_1118_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1724_ ) );
OAI21_X1 \myreg/_4211_ ( .A(\myreg/_1724_ ), .B1(\myreg/_0122_ ), .B2(fanout_net_46 ), .ZN(\myreg/_1725_ ) );
AOI21_X1 \myreg/_4212_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1723_ ), .B2(\myreg/_1725_ ), .ZN(\myreg/_1726_ ) );
OR2_X1 \myreg/_4213_ ( .A1(\myreg/_1721_ ), .A2(\myreg/_1726_ ), .ZN(\myreg/_1727_ ) );
MUX2_X1 \myreg/_4214_ ( .A(\myreg/_0346_ ), .B(\myreg/_0378_ ), .S(fanout_net_46 ), .Z(\myreg/_1728_ ) );
MUX2_X1 \myreg/_4215_ ( .A(\myreg/_0410_ ), .B(\myreg/_0442_ ), .S(fanout_net_46 ), .Z(\myreg/_1729_ ) );
MUX2_X1 \myreg/_4216_ ( .A(\myreg/_1728_ ), .B(\myreg/_1729_ ), .S(fanout_net_54 ), .Z(\myreg/_1730_ ) );
MUX2_X1 \myreg/_4217_ ( .A(\myreg/_0026_ ), .B(\myreg/_0250_ ), .S(fanout_net_46 ), .Z(\myreg/_1731_ ) );
MUX2_X1 \myreg/_4218_ ( .A(\myreg/_0282_ ), .B(\myreg/_0314_ ), .S(fanout_net_46 ), .Z(\myreg/_1732_ ) );
MUX2_X1 \myreg/_4219_ ( .A(\myreg/_1731_ ), .B(\myreg/_1732_ ), .S(fanout_net_54 ), .Z(\myreg/_1733_ ) );
MUX2_X1 \myreg/_4220_ ( .A(\myreg/_1730_ ), .B(\myreg/_1733_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1734_ ) );
MUX2_X1 \myreg/_4221_ ( .A(\myreg/_1727_ ), .B(\myreg/_1734_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2406_ ) );
MUX2_X1 \myreg/_4222_ ( .A(\myreg/_0475_ ), .B(\myreg/_0507_ ), .S(fanout_net_46 ), .Z(\myreg/_1735_ ) );
MUX2_X1 \myreg/_4223_ ( .A(\myreg/_0059_ ), .B(\myreg/_0091_ ), .S(fanout_net_46 ), .Z(\myreg/_1736_ ) );
MUX2_X1 \myreg/_4224_ ( .A(\myreg/_1735_ ), .B(\myreg/_1736_ ), .S(fanout_net_55 ), .Z(\myreg/_1737_ ) );
MUX2_X1 \myreg/_4225_ ( .A(\myreg/_0123_ ), .B(\myreg/_0155_ ), .S(fanout_net_46 ), .Z(\myreg/_1738_ ) );
MUX2_X1 \myreg/_4226_ ( .A(\myreg/_0187_ ), .B(\myreg/_0219_ ), .S(fanout_net_46 ), .Z(\myreg/_1739_ ) );
MUX2_X1 \myreg/_4227_ ( .A(\myreg/_1738_ ), .B(\myreg/_1739_ ), .S(fanout_net_55 ), .Z(\myreg/_1740_ ) );
MUX2_X1 \myreg/_4228_ ( .A(\myreg/_1737_ ), .B(\myreg/_1740_ ), .S(fanout_net_60 ), .Z(\myreg/_1741_ ) );
MUX2_X1 \myreg/_4229_ ( .A(\myreg/_0347_ ), .B(\myreg/_0379_ ), .S(fanout_net_46 ), .Z(\myreg/_1742_ ) );
MUX2_X1 \myreg/_4230_ ( .A(\myreg/_0411_ ), .B(\myreg/_0443_ ), .S(fanout_net_46 ), .Z(\myreg/_1743_ ) );
MUX2_X1 \myreg/_4231_ ( .A(\myreg/_1742_ ), .B(\myreg/_1743_ ), .S(fanout_net_55 ), .Z(\myreg/_1744_ ) );
MUX2_X1 \myreg/_4232_ ( .A(\myreg/_0027_ ), .B(\myreg/_0251_ ), .S(fanout_net_46 ), .Z(\myreg/_1745_ ) );
MUX2_X1 \myreg/_4233_ ( .A(\myreg/_0283_ ), .B(\myreg/_0315_ ), .S(fanout_net_46 ), .Z(\myreg/_1746_ ) );
MUX2_X1 \myreg/_4234_ ( .A(\myreg/_1745_ ), .B(\myreg/_1746_ ), .S(fanout_net_55 ), .Z(\myreg/_1747_ ) );
MUX2_X1 \myreg/_4235_ ( .A(\myreg/_1744_ ), .B(\myreg/_1747_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1748_ ) );
MUX2_X1 \myreg/_4236_ ( .A(\myreg/_1741_ ), .B(\myreg/_1748_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2407_ ) );
MUX2_X1 \myreg/_4237_ ( .A(\myreg/_0476_ ), .B(\myreg/_0508_ ), .S(fanout_net_46 ), .Z(\myreg/_1749_ ) );
MUX2_X1 \myreg/_4238_ ( .A(\myreg/_0060_ ), .B(\myreg/_0092_ ), .S(fanout_net_47 ), .Z(\myreg/_1750_ ) );
MUX2_X1 \myreg/_4239_ ( .A(\myreg/_1749_ ), .B(\myreg/_1750_ ), .S(fanout_net_55 ), .Z(\myreg/_1751_ ) );
MUX2_X1 \myreg/_4240_ ( .A(\myreg/_0124_ ), .B(\myreg/_0156_ ), .S(fanout_net_47 ), .Z(\myreg/_1752_ ) );
MUX2_X1 \myreg/_4241_ ( .A(\myreg/_0188_ ), .B(\myreg/_0220_ ), .S(fanout_net_47 ), .Z(\myreg/_1753_ ) );
MUX2_X1 \myreg/_4242_ ( .A(\myreg/_1752_ ), .B(\myreg/_1753_ ), .S(fanout_net_55 ), .Z(\myreg/_1754_ ) );
MUX2_X1 \myreg/_4243_ ( .A(\myreg/_1751_ ), .B(\myreg/_1754_ ), .S(fanout_net_60 ), .Z(\myreg/_1755_ ) );
MUX2_X1 \myreg/_4244_ ( .A(\myreg/_0348_ ), .B(\myreg/_0380_ ), .S(fanout_net_47 ), .Z(\myreg/_1756_ ) );
MUX2_X1 \myreg/_4245_ ( .A(\myreg/_0412_ ), .B(\myreg/_0444_ ), .S(fanout_net_47 ), .Z(\myreg/_1757_ ) );
MUX2_X1 \myreg/_4246_ ( .A(\myreg/_1756_ ), .B(\myreg/_1757_ ), .S(fanout_net_55 ), .Z(\myreg/_1758_ ) );
MUX2_X1 \myreg/_4247_ ( .A(\myreg/_0028_ ), .B(\myreg/_0252_ ), .S(fanout_net_47 ), .Z(\myreg/_1759_ ) );
MUX2_X1 \myreg/_4248_ ( .A(\myreg/_0284_ ), .B(\myreg/_0316_ ), .S(fanout_net_47 ), .Z(\myreg/_1760_ ) );
MUX2_X1 \myreg/_4249_ ( .A(\myreg/_1759_ ), .B(\myreg/_1760_ ), .S(fanout_net_55 ), .Z(\myreg/_1761_ ) );
MUX2_X1 \myreg/_4250_ ( .A(\myreg/_1758_ ), .B(\myreg/_1761_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1762_ ) );
MUX2_X1 \myreg/_4251_ ( .A(\myreg/_1755_ ), .B(\myreg/_1762_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2408_ ) );
MUX2_X1 \myreg/_4252_ ( .A(\myreg/_0477_ ), .B(\myreg/_0509_ ), .S(fanout_net_47 ), .Z(\myreg/_1763_ ) );
MUX2_X1 \myreg/_4253_ ( .A(\myreg/_0061_ ), .B(\myreg/_0093_ ), .S(fanout_net_47 ), .Z(\myreg/_1764_ ) );
MUX2_X1 \myreg/_4254_ ( .A(\myreg/_1763_ ), .B(\myreg/_1764_ ), .S(fanout_net_55 ), .Z(\myreg/_1765_ ) );
MUX2_X1 \myreg/_4255_ ( .A(\myreg/_0125_ ), .B(\myreg/_0157_ ), .S(fanout_net_47 ), .Z(\myreg/_1766_ ) );
MUX2_X1 \myreg/_4256_ ( .A(\myreg/_0189_ ), .B(\myreg/_0221_ ), .S(fanout_net_47 ), .Z(\myreg/_1767_ ) );
MUX2_X1 \myreg/_4257_ ( .A(\myreg/_1766_ ), .B(\myreg/_1767_ ), .S(fanout_net_55 ), .Z(\myreg/_1768_ ) );
MUX2_X1 \myreg/_4258_ ( .A(\myreg/_1765_ ), .B(\myreg/_1768_ ), .S(fanout_net_60 ), .Z(\myreg/_1769_ ) );
MUX2_X1 \myreg/_4259_ ( .A(\myreg/_0349_ ), .B(\myreg/_0381_ ), .S(fanout_net_47 ), .Z(\myreg/_1770_ ) );
MUX2_X1 \myreg/_4260_ ( .A(\myreg/_0413_ ), .B(\myreg/_0445_ ), .S(fanout_net_47 ), .Z(\myreg/_1771_ ) );
MUX2_X1 \myreg/_4261_ ( .A(\myreg/_1770_ ), .B(\myreg/_1771_ ), .S(fanout_net_55 ), .Z(\myreg/_1772_ ) );
MUX2_X1 \myreg/_4262_ ( .A(\myreg/_0029_ ), .B(\myreg/_0253_ ), .S(fanout_net_47 ), .Z(\myreg/_1773_ ) );
MUX2_X1 \myreg/_4263_ ( .A(\myreg/_0285_ ), .B(\myreg/_0317_ ), .S(fanout_net_47 ), .Z(\myreg/_1774_ ) );
MUX2_X1 \myreg/_4264_ ( .A(\myreg/_1773_ ), .B(\myreg/_1774_ ), .S(fanout_net_55 ), .Z(\myreg/_1775_ ) );
MUX2_X1 \myreg/_4265_ ( .A(\myreg/_1772_ ), .B(\myreg/_1775_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1776_ ) );
MUX2_X1 \myreg/_4266_ ( .A(\myreg/_1769_ ), .B(\myreg/_1776_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2409_ ) );
OR2_X1 \myreg/_4267_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0222_ ), .ZN(\myreg/_1777_ ) );
OAI211_X2 \myreg/_4268_ ( .A(\myreg/_1777_ ), .B(fanout_net_55 ), .C1(\myreg/_0190_ ), .C2(fanout_net_47 ), .ZN(\myreg/_1778_ ) );
AOI21_X1 \myreg/_4269_ ( .A(fanout_net_55 ), .B1(\myreg/_1181_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1779_ ) );
OAI21_X1 \myreg/_4270_ ( .A(\myreg/_1779_ ), .B1(\myreg/_0126_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1780_ ) );
AOI21_X1 \myreg/_4271_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1778_ ), .B2(\myreg/_1780_ ), .ZN(\myreg/_1781_ ) );
OR2_X1 \myreg/_4272_ ( .A1(\myreg/_0062_ ), .A2(fanout_net_47 ), .ZN(\myreg/_1782_ ) );
OAI211_X2 \myreg/_4273_ ( .A(\myreg/_1782_ ), .B(fanout_net_55 ), .C1(\myreg/_0094_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1783_ ) );
AOI21_X1 \myreg/_4274_ ( .A(fanout_net_55 ), .B1(\myreg/_1187_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1784_ ) );
OAI21_X1 \myreg/_4275_ ( .A(\myreg/_1784_ ), .B1(\myreg/_0478_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1785_ ) );
AOI21_X1 \myreg/_4276_ ( .A(fanout_net_60 ), .B1(\myreg/_1783_ ), .B2(\myreg/_1785_ ), .ZN(\myreg/_1786_ ) );
OR2_X1 \myreg/_4277_ ( .A1(\myreg/_1781_ ), .A2(\myreg/_1786_ ), .ZN(\myreg/_1787_ ) );
MUX2_X1 \myreg/_4278_ ( .A(\myreg/_0350_ ), .B(\myreg/_0382_ ), .S(fanout_net_47 ), .Z(\myreg/_1788_ ) );
MUX2_X1 \myreg/_4279_ ( .A(\myreg/_0414_ ), .B(\myreg/_0446_ ), .S(fanout_net_47 ), .Z(\myreg/_1789_ ) );
MUX2_X1 \myreg/_4280_ ( .A(\myreg/_1788_ ), .B(\myreg/_1789_ ), .S(fanout_net_55 ), .Z(\myreg/_1790_ ) );
MUX2_X1 \myreg/_4281_ ( .A(\myreg/_0030_ ), .B(\myreg/_0254_ ), .S(fanout_net_47 ), .Z(\myreg/_1791_ ) );
MUX2_X1 \myreg/_4282_ ( .A(\myreg/_0286_ ), .B(\myreg/_0318_ ), .S(fanout_net_47 ), .Z(\myreg/_1792_ ) );
MUX2_X1 \myreg/_4283_ ( .A(\myreg/_1791_ ), .B(\myreg/_1792_ ), .S(fanout_net_55 ), .Z(\myreg/_1793_ ) );
MUX2_X1 \myreg/_4284_ ( .A(\myreg/_1790_ ), .B(\myreg/_1793_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1794_ ) );
MUX2_X1 \myreg/_4285_ ( .A(\myreg/_1787_ ), .B(\myreg/_1794_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2410_ ) );
OR2_X1 \myreg/_4286_ ( .A1(\myreg/_1679_ ), .A2(\myreg/_0223_ ), .ZN(\myreg/_1795_ ) );
OAI211_X2 \myreg/_4287_ ( .A(\myreg/_1795_ ), .B(fanout_net_55 ), .C1(\myreg/_0191_ ), .C2(fanout_net_47 ), .ZN(\myreg/_1796_ ) );
AOI21_X1 \myreg/_4288_ ( .A(fanout_net_55 ), .B1(\myreg/_1208_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1797_ ) );
OAI21_X1 \myreg/_4289_ ( .A(\myreg/_1797_ ), .B1(\myreg/_0127_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1798_ ) );
NAND3_X1 \myreg/_4290_ ( .A1(\myreg/_1796_ ), .A2(fanout_net_60 ), .A3(\myreg/_1798_ ), .ZN(\myreg/_1799_ ) );
OR2_X1 \myreg/_4291_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0095_ ), .ZN(\myreg/_1800_ ) );
OAI211_X2 \myreg/_4292_ ( .A(\myreg/_1800_ ), .B(fanout_net_55 ), .C1(\myreg/_0063_ ), .C2(fanout_net_47 ), .ZN(\myreg/_1801_ ) );
AOI21_X1 \myreg/_4293_ ( .A(fanout_net_55 ), .B1(\myreg/_1202_ ), .B2(fanout_net_47 ), .ZN(\myreg/_1802_ ) );
OAI21_X1 \myreg/_4294_ ( .A(\myreg/_1802_ ), .B1(\myreg/_0479_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1803_ ) );
NAND3_X1 \myreg/_4295_ ( .A1(\myreg/_1801_ ), .A2(\myreg/_1656_ ), .A3(\myreg/_1803_ ), .ZN(\myreg/_1804_ ) );
AND2_X1 \myreg/_4296_ ( .A1(\myreg/_1799_ ), .A2(\myreg/_1804_ ), .ZN(\myreg/_1805_ ) );
MUX2_X1 \myreg/_4297_ ( .A(\myreg/_0351_ ), .B(\myreg/_0383_ ), .S(fanout_net_48 ), .Z(\myreg/_1806_ ) );
MUX2_X1 \myreg/_4298_ ( .A(\myreg/_0415_ ), .B(\myreg/_0447_ ), .S(fanout_net_48 ), .Z(\myreg/_1807_ ) );
MUX2_X1 \myreg/_4299_ ( .A(\myreg/_1806_ ), .B(\myreg/_1807_ ), .S(fanout_net_55 ), .Z(\myreg/_1808_ ) );
MUX2_X1 \myreg/_4300_ ( .A(\myreg/_0031_ ), .B(\myreg/_0255_ ), .S(fanout_net_48 ), .Z(\myreg/_1809_ ) );
MUX2_X1 \myreg/_4301_ ( .A(\myreg/_0287_ ), .B(\myreg/_0319_ ), .S(fanout_net_48 ), .Z(\myreg/_1810_ ) );
MUX2_X1 \myreg/_4302_ ( .A(\myreg/_1809_ ), .B(\myreg/_1810_ ), .S(fanout_net_55 ), .Z(\myreg/_1811_ ) );
MUX2_X1 \myreg/_4303_ ( .A(\myreg/_1808_ ), .B(\myreg/_1811_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1812_ ) );
MUX2_X1 \myreg/_4304_ ( .A(\myreg/_1805_ ), .B(\myreg/_1812_ ), .S(\myreg/_1659_ ), .Z(\myreg/_2411_ ) );
OR2_X1 \myreg/_4305_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0193_ ), .ZN(\myreg/_1813_ ) );
OAI211_X2 \myreg/_4306_ ( .A(\myreg/_1813_ ), .B(fanout_net_55 ), .C1(\myreg/_0161_ ), .C2(fanout_net_48 ), .ZN(\myreg/_1814_ ) );
AOI21_X1 \myreg/_4307_ ( .A(fanout_net_55 ), .B1(\myreg/_1222_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1815_ ) );
OAI21_X1 \myreg/_4308_ ( .A(\myreg/_1815_ ), .B1(\myreg/_0097_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1816_ ) );
AOI21_X1 \myreg/_4309_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1814_ ), .B2(\myreg/_1816_ ), .ZN(\myreg/_1817_ ) );
OR2_X1 \myreg/_4310_ ( .A1(\myreg/_0033_ ), .A2(fanout_net_48 ), .ZN(\myreg/_1818_ ) );
OAI211_X2 \myreg/_4311_ ( .A(\myreg/_1818_ ), .B(fanout_net_55 ), .C1(\myreg/_0065_ ), .C2(\myreg/_1679_ ), .ZN(\myreg/_1819_ ) );
AOI21_X1 \myreg/_4312_ ( .A(fanout_net_55 ), .B1(\myreg/_1229_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1820_ ) );
OAI21_X1 \myreg/_4313_ ( .A(\myreg/_1820_ ), .B1(\myreg/_0449_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1821_ ) );
AOI21_X1 \myreg/_4314_ ( .A(fanout_net_60 ), .B1(\myreg/_1819_ ), .B2(\myreg/_1821_ ), .ZN(\myreg/_1822_ ) );
OR2_X1 \myreg/_4315_ ( .A1(\myreg/_1817_ ), .A2(\myreg/_1822_ ), .ZN(\myreg/_1823_ ) );
MUX2_X1 \myreg/_4316_ ( .A(\myreg/_0321_ ), .B(\myreg/_0353_ ), .S(fanout_net_48 ), .Z(\myreg/_1824_ ) );
MUX2_X1 \myreg/_4317_ ( .A(\myreg/_0385_ ), .B(\myreg/_0417_ ), .S(fanout_net_48 ), .Z(\myreg/_1825_ ) );
MUX2_X1 \myreg/_4318_ ( .A(\myreg/_1824_ ), .B(\myreg/_1825_ ), .S(fanout_net_55 ), .Z(\myreg/_1826_ ) );
MUX2_X1 \myreg/_4319_ ( .A(\myreg/_0001_ ), .B(\myreg/_0225_ ), .S(fanout_net_48 ), .Z(\myreg/_1827_ ) );
MUX2_X1 \myreg/_4320_ ( .A(\myreg/_0257_ ), .B(\myreg/_0289_ ), .S(fanout_net_48 ), .Z(\myreg/_1828_ ) );
MUX2_X1 \myreg/_4321_ ( .A(\myreg/_1827_ ), .B(\myreg/_1828_ ), .S(fanout_net_55 ), .Z(\myreg/_1829_ ) );
MUX2_X1 \myreg/_4322_ ( .A(\myreg/_1826_ ), .B(\myreg/_1829_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1830_ ) );
BUF_X4 \myreg/_4323_ ( .A(\myreg/_1658_ ), .Z(\myreg/_1831_ ) );
MUX2_X1 \myreg/_4324_ ( .A(\myreg/_1823_ ), .B(\myreg/_1830_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2381_ ) );
MUX2_X1 \myreg/_4325_ ( .A(\myreg/_0450_ ), .B(\myreg/_0482_ ), .S(fanout_net_48 ), .Z(\myreg/_1832_ ) );
MUX2_X1 \myreg/_4326_ ( .A(\myreg/_0034_ ), .B(\myreg/_0066_ ), .S(fanout_net_48 ), .Z(\myreg/_1833_ ) );
MUX2_X1 \myreg/_4327_ ( .A(\myreg/_1832_ ), .B(\myreg/_1833_ ), .S(fanout_net_56 ), .Z(\myreg/_1834_ ) );
MUX2_X1 \myreg/_4328_ ( .A(\myreg/_0098_ ), .B(\myreg/_0130_ ), .S(fanout_net_48 ), .Z(\myreg/_1835_ ) );
MUX2_X1 \myreg/_4329_ ( .A(\myreg/_0162_ ), .B(\myreg/_0194_ ), .S(fanout_net_48 ), .Z(\myreg/_1836_ ) );
MUX2_X1 \myreg/_4330_ ( .A(\myreg/_1835_ ), .B(\myreg/_1836_ ), .S(fanout_net_56 ), .Z(\myreg/_1837_ ) );
MUX2_X1 \myreg/_4331_ ( .A(\myreg/_1834_ ), .B(\myreg/_1837_ ), .S(fanout_net_60 ), .Z(\myreg/_1838_ ) );
MUX2_X1 \myreg/_4332_ ( .A(\myreg/_0322_ ), .B(\myreg/_0354_ ), .S(fanout_net_48 ), .Z(\myreg/_1839_ ) );
MUX2_X1 \myreg/_4333_ ( .A(\myreg/_0386_ ), .B(\myreg/_0418_ ), .S(fanout_net_48 ), .Z(\myreg/_1840_ ) );
MUX2_X1 \myreg/_4334_ ( .A(\myreg/_1839_ ), .B(\myreg/_1840_ ), .S(fanout_net_56 ), .Z(\myreg/_1841_ ) );
MUX2_X1 \myreg/_4335_ ( .A(\myreg/_0002_ ), .B(\myreg/_0226_ ), .S(fanout_net_48 ), .Z(\myreg/_1842_ ) );
MUX2_X1 \myreg/_4336_ ( .A(\myreg/_0258_ ), .B(\myreg/_0290_ ), .S(fanout_net_48 ), .Z(\myreg/_1843_ ) );
MUX2_X1 \myreg/_4337_ ( .A(\myreg/_1842_ ), .B(\myreg/_1843_ ), .S(fanout_net_56 ), .Z(\myreg/_1844_ ) );
MUX2_X1 \myreg/_4338_ ( .A(\myreg/_1841_ ), .B(\myreg/_1844_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1845_ ) );
MUX2_X1 \myreg/_4339_ ( .A(\myreg/_1838_ ), .B(\myreg/_1845_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2382_ ) );
OR2_X1 \myreg/_4340_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0067_ ), .ZN(\myreg/_1846_ ) );
OAI211_X2 \myreg/_4341_ ( .A(\myreg/_1846_ ), .B(fanout_net_56 ), .C1(\myreg/_0035_ ), .C2(fanout_net_48 ), .ZN(\myreg/_1847_ ) );
AOI21_X1 \myreg/_4342_ ( .A(fanout_net_56 ), .B1(\myreg/_1258_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1848_ ) );
OAI21_X1 \myreg/_4343_ ( .A(\myreg/_1848_ ), .B1(\myreg/_0451_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1849_ ) );
AOI21_X1 \myreg/_4344_ ( .A(fanout_net_60 ), .B1(\myreg/_1847_ ), .B2(\myreg/_1849_ ), .ZN(\myreg/_1850_ ) );
OR2_X1 \myreg/_4345_ ( .A1(\myreg/_0163_ ), .A2(fanout_net_48 ), .ZN(\myreg/_1851_ ) );
OAI211_X2 \myreg/_4346_ ( .A(\myreg/_1851_ ), .B(fanout_net_56 ), .C1(\myreg/_0195_ ), .C2(\myreg/_1679_ ), .ZN(\myreg/_1852_ ) );
AOI21_X1 \myreg/_4347_ ( .A(fanout_net_56 ), .B1(\myreg/_1264_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1853_ ) );
OAI21_X1 \myreg/_4348_ ( .A(\myreg/_1853_ ), .B1(\myreg/_0099_ ), .B2(fanout_net_48 ), .ZN(\myreg/_1854_ ) );
AOI21_X1 \myreg/_4349_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1852_ ), .B2(\myreg/_1854_ ), .ZN(\myreg/_1855_ ) );
OR2_X1 \myreg/_4350_ ( .A1(\myreg/_1850_ ), .A2(\myreg/_1855_ ), .ZN(\myreg/_1856_ ) );
MUX2_X1 \myreg/_4351_ ( .A(\myreg/_0323_ ), .B(\myreg/_0355_ ), .S(fanout_net_48 ), .Z(\myreg/_1857_ ) );
MUX2_X1 \myreg/_4352_ ( .A(\myreg/_0387_ ), .B(\myreg/_0419_ ), .S(fanout_net_49 ), .Z(\myreg/_1858_ ) );
MUX2_X1 \myreg/_4353_ ( .A(\myreg/_1857_ ), .B(\myreg/_1858_ ), .S(fanout_net_56 ), .Z(\myreg/_1859_ ) );
MUX2_X1 \myreg/_4354_ ( .A(\myreg/_0003_ ), .B(\myreg/_0227_ ), .S(fanout_net_49 ), .Z(\myreg/_1860_ ) );
MUX2_X1 \myreg/_4355_ ( .A(\myreg/_0259_ ), .B(\myreg/_0291_ ), .S(fanout_net_49 ), .Z(\myreg/_1861_ ) );
MUX2_X1 \myreg/_4356_ ( .A(\myreg/_1860_ ), .B(\myreg/_1861_ ), .S(fanout_net_56 ), .Z(\myreg/_1862_ ) );
MUX2_X1 \myreg/_4357_ ( .A(\myreg/_1859_ ), .B(\myreg/_1862_ ), .S(\myreg/_1715_ ), .Z(\myreg/_1863_ ) );
MUX2_X1 \myreg/_4358_ ( .A(\myreg/_1856_ ), .B(\myreg/_1863_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2383_ ) );
MUX2_X1 \myreg/_4359_ ( .A(\myreg/_0100_ ), .B(\myreg/_0132_ ), .S(fanout_net_49 ), .Z(\myreg/_1864_ ) );
MUX2_X1 \myreg/_4360_ ( .A(\myreg/_0164_ ), .B(\myreg/_0196_ ), .S(fanout_net_49 ), .Z(\myreg/_1865_ ) );
MUX2_X1 \myreg/_4361_ ( .A(\myreg/_1864_ ), .B(\myreg/_1865_ ), .S(fanout_net_56 ), .Z(\myreg/_1866_ ) );
MUX2_X1 \myreg/_4362_ ( .A(\myreg/_0452_ ), .B(\myreg/_0484_ ), .S(fanout_net_49 ), .Z(\myreg/_1867_ ) );
MUX2_X1 \myreg/_4363_ ( .A(\myreg/_0036_ ), .B(\myreg/_0068_ ), .S(fanout_net_49 ), .Z(\myreg/_1868_ ) );
MUX2_X1 \myreg/_4364_ ( .A(\myreg/_1867_ ), .B(\myreg/_1868_ ), .S(fanout_net_56 ), .Z(\myreg/_1869_ ) );
MUX2_X1 \myreg/_4365_ ( .A(\myreg/_1866_ ), .B(\myreg/_1869_ ), .S(\myreg/_1660_ ), .Z(\myreg/_1870_ ) );
MUX2_X1 \myreg/_4366_ ( .A(\myreg/_0004_ ), .B(\myreg/_0260_ ), .S(fanout_net_56 ), .Z(\myreg/_1871_ ) );
MUX2_X1 \myreg/_4367_ ( .A(\myreg/_0228_ ), .B(\myreg/_0292_ ), .S(fanout_net_56 ), .Z(\myreg/_1872_ ) );
MUX2_X1 \myreg/_4368_ ( .A(\myreg/_1871_ ), .B(\myreg/_1872_ ), .S(fanout_net_49 ), .Z(\myreg/_1873_ ) );
MUX2_X1 \myreg/_4369_ ( .A(\myreg/_0324_ ), .B(\myreg/_0388_ ), .S(fanout_net_56 ), .Z(\myreg/_1874_ ) );
MUX2_X1 \myreg/_4370_ ( .A(\myreg/_0356_ ), .B(\myreg/_0420_ ), .S(fanout_net_56 ), .Z(\myreg/_1875_ ) );
MUX2_X1 \myreg/_4371_ ( .A(\myreg/_1874_ ), .B(\myreg/_1875_ ), .S(fanout_net_49 ), .Z(\myreg/_1876_ ) );
MUX2_X1 \myreg/_4372_ ( .A(\myreg/_1873_ ), .B(\myreg/_1876_ ), .S(fanout_net_60 ), .Z(\myreg/_1877_ ) );
MUX2_X1 \myreg/_4373_ ( .A(\myreg/_1870_ ), .B(\myreg/_1877_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2384_ ) );
OR2_X1 \myreg/_4374_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0197_ ), .ZN(\myreg/_1878_ ) );
OAI211_X2 \myreg/_4375_ ( .A(\myreg/_1878_ ), .B(fanout_net_56 ), .C1(\myreg/_0165_ ), .C2(fanout_net_49 ), .ZN(\myreg/_1879_ ) );
AOI21_X1 \myreg/_4376_ ( .A(fanout_net_56 ), .B1(\myreg/_1304_ ), .B2(fanout_net_49 ), .ZN(\myreg/_1880_ ) );
OAI21_X1 \myreg/_4377_ ( .A(\myreg/_1880_ ), .B1(\myreg/_0101_ ), .B2(fanout_net_49 ), .ZN(\myreg/_1881_ ) );
AOI21_X1 \myreg/_4378_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1879_ ), .B2(\myreg/_1881_ ), .ZN(\myreg/_1882_ ) );
OR2_X1 \myreg/_4379_ ( .A1(\myreg/_0037_ ), .A2(fanout_net_49 ), .ZN(\myreg/_1883_ ) );
OAI211_X2 \myreg/_4380_ ( .A(\myreg/_1883_ ), .B(fanout_net_56 ), .C1(\myreg/_0069_ ), .C2(\myreg/_1679_ ), .ZN(\myreg/_1884_ ) );
AOI21_X1 \myreg/_4381_ ( .A(fanout_net_56 ), .B1(\myreg/_1298_ ), .B2(fanout_net_49 ), .ZN(\myreg/_1885_ ) );
OAI21_X1 \myreg/_4382_ ( .A(\myreg/_1885_ ), .B1(\myreg/_0453_ ), .B2(fanout_net_49 ), .ZN(\myreg/_1886_ ) );
AOI21_X1 \myreg/_4383_ ( .A(fanout_net_60 ), .B1(\myreg/_1884_ ), .B2(\myreg/_1886_ ), .ZN(\myreg/_1887_ ) );
OR2_X1 \myreg/_4384_ ( .A1(\myreg/_1882_ ), .A2(\myreg/_1887_ ), .ZN(\myreg/_1888_ ) );
MUX2_X1 \myreg/_4385_ ( .A(\myreg/_0325_ ), .B(\myreg/_0357_ ), .S(fanout_net_49 ), .Z(\myreg/_1889_ ) );
MUX2_X1 \myreg/_4386_ ( .A(\myreg/_0389_ ), .B(\myreg/_0421_ ), .S(fanout_net_49 ), .Z(\myreg/_1890_ ) );
MUX2_X1 \myreg/_4387_ ( .A(\myreg/_1889_ ), .B(\myreg/_1890_ ), .S(fanout_net_56 ), .Z(\myreg/_1891_ ) );
MUX2_X1 \myreg/_4388_ ( .A(\myreg/_0005_ ), .B(\myreg/_0229_ ), .S(fanout_net_49 ), .Z(\myreg/_1892_ ) );
MUX2_X1 \myreg/_4389_ ( .A(\myreg/_0261_ ), .B(\myreg/_0293_ ), .S(fanout_net_49 ), .Z(\myreg/_1893_ ) );
MUX2_X1 \myreg/_4390_ ( .A(\myreg/_1892_ ), .B(\myreg/_1893_ ), .S(fanout_net_56 ), .Z(\myreg/_1894_ ) );
BUF_X4 \myreg/_4391_ ( .A(\myreg/_1641_ ), .Z(\myreg/_1895_ ) );
MUX2_X1 \myreg/_4392_ ( .A(\myreg/_1891_ ), .B(\myreg/_1894_ ), .S(\myreg/_1895_ ), .Z(\myreg/_1896_ ) );
MUX2_X1 \myreg/_4393_ ( .A(\myreg/_1888_ ), .B(\myreg/_1896_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2385_ ) );
MUX2_X1 \myreg/_4394_ ( .A(\myreg/_0454_ ), .B(\myreg/_0486_ ), .S(fanout_net_49 ), .Z(\myreg/_1897_ ) );
MUX2_X1 \myreg/_4395_ ( .A(\myreg/_0038_ ), .B(\myreg/_0070_ ), .S(fanout_net_49 ), .Z(\myreg/_1898_ ) );
MUX2_X1 \myreg/_4396_ ( .A(\myreg/_1897_ ), .B(\myreg/_1898_ ), .S(fanout_net_56 ), .Z(\myreg/_1899_ ) );
MUX2_X1 \myreg/_4397_ ( .A(\myreg/_0102_ ), .B(\myreg/_0134_ ), .S(fanout_net_49 ), .Z(\myreg/_1900_ ) );
MUX2_X1 \myreg/_4398_ ( .A(\myreg/_0166_ ), .B(\myreg/_0198_ ), .S(fanout_net_49 ), .Z(\myreg/_1901_ ) );
MUX2_X1 \myreg/_4399_ ( .A(\myreg/_1900_ ), .B(\myreg/_1901_ ), .S(fanout_net_56 ), .Z(\myreg/_1902_ ) );
MUX2_X1 \myreg/_4400_ ( .A(\myreg/_1899_ ), .B(\myreg/_1902_ ), .S(fanout_net_60 ), .Z(\myreg/_1903_ ) );
MUX2_X1 \myreg/_4401_ ( .A(\myreg/_0326_ ), .B(\myreg/_0358_ ), .S(fanout_net_49 ), .Z(\myreg/_1904_ ) );
MUX2_X1 \myreg/_4402_ ( .A(\myreg/_0390_ ), .B(\myreg/_0422_ ), .S(fanout_net_49 ), .Z(\myreg/_1905_ ) );
MUX2_X1 \myreg/_4403_ ( .A(\myreg/_1904_ ), .B(\myreg/_1905_ ), .S(fanout_net_56 ), .Z(\myreg/_1906_ ) );
MUX2_X1 \myreg/_4404_ ( .A(\myreg/_0006_ ), .B(\myreg/_0230_ ), .S(fanout_net_49 ), .Z(\myreg/_1907_ ) );
MUX2_X1 \myreg/_4405_ ( .A(\myreg/_0262_ ), .B(\myreg/_0294_ ), .S(fanout_net_49 ), .Z(\myreg/_1908_ ) );
MUX2_X1 \myreg/_4406_ ( .A(\myreg/_1907_ ), .B(\myreg/_1908_ ), .S(fanout_net_56 ), .Z(\myreg/_1909_ ) );
MUX2_X1 \myreg/_4407_ ( .A(\myreg/_1906_ ), .B(\myreg/_1909_ ), .S(\myreg/_1895_ ), .Z(\myreg/_1910_ ) );
MUX2_X1 \myreg/_4408_ ( .A(\myreg/_1903_ ), .B(\myreg/_1910_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2386_ ) );
OR2_X1 \myreg/_4409_ ( .A1(\myreg/_0167_ ), .A2(fanout_net_49 ), .ZN(\myreg/_1911_ ) );
OAI211_X2 \myreg/_4410_ ( .A(\myreg/_1911_ ), .B(fanout_net_56 ), .C1(\myreg/_0199_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1912_ ) );
AOI21_X1 \myreg/_4411_ ( .A(fanout_net_56 ), .B1(\myreg/_1332_ ), .B2(fanout_net_49 ), .ZN(\myreg/_1913_ ) );
OAI21_X1 \myreg/_4412_ ( .A(\myreg/_1913_ ), .B1(\myreg/_0103_ ), .B2(fanout_net_49 ), .ZN(\myreg/_1914_ ) );
NAND3_X1 \myreg/_4413_ ( .A1(\myreg/_1912_ ), .A2(\myreg/_1914_ ), .A3(fanout_net_60 ), .ZN(\myreg/_1915_ ) );
OR2_X1 \myreg/_4414_ ( .A1(\myreg/_0039_ ), .A2(fanout_net_50 ), .ZN(\myreg/_1916_ ) );
OAI211_X2 \myreg/_4415_ ( .A(\myreg/_1916_ ), .B(fanout_net_56 ), .C1(\myreg/_0071_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_1917_ ) );
AOI21_X1 \myreg/_4416_ ( .A(fanout_net_56 ), .B1(\myreg/_1338_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1918_ ) );
OAI21_X1 \myreg/_4417_ ( .A(\myreg/_1918_ ), .B1(\myreg/_0455_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1919_ ) );
NAND3_X1 \myreg/_4418_ ( .A1(\myreg/_1917_ ), .A2(\myreg/_1919_ ), .A3(\myreg/_1656_ ), .ZN(\myreg/_1920_ ) );
AND2_X1 \myreg/_4419_ ( .A1(\myreg/_1915_ ), .A2(\myreg/_1920_ ), .ZN(\myreg/_1921_ ) );
MUX2_X1 \myreg/_4420_ ( .A(\myreg/_0327_ ), .B(\myreg/_0359_ ), .S(fanout_net_50 ), .Z(\myreg/_1922_ ) );
MUX2_X1 \myreg/_4421_ ( .A(\myreg/_0391_ ), .B(\myreg/_0423_ ), .S(fanout_net_50 ), .Z(\myreg/_1923_ ) );
MUX2_X1 \myreg/_4422_ ( .A(\myreg/_1922_ ), .B(\myreg/_1923_ ), .S(fanout_net_57 ), .Z(\myreg/_1924_ ) );
MUX2_X1 \myreg/_4423_ ( .A(\myreg/_0007_ ), .B(\myreg/_0231_ ), .S(fanout_net_50 ), .Z(\myreg/_1925_ ) );
MUX2_X1 \myreg/_4424_ ( .A(\myreg/_0263_ ), .B(\myreg/_0295_ ), .S(fanout_net_50 ), .Z(\myreg/_1926_ ) );
MUX2_X1 \myreg/_4425_ ( .A(\myreg/_1925_ ), .B(\myreg/_1926_ ), .S(fanout_net_57 ), .Z(\myreg/_1927_ ) );
MUX2_X1 \myreg/_4426_ ( .A(\myreg/_1924_ ), .B(\myreg/_1927_ ), .S(\myreg/_1895_ ), .Z(\myreg/_1928_ ) );
MUX2_X1 \myreg/_4427_ ( .A(\myreg/_1921_ ), .B(\myreg/_1928_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2387_ ) );
OR2_X1 \myreg/_4428_ ( .A1(\myreg/_1634_ ), .A2(\myreg/_0200_ ), .ZN(\myreg/_1929_ ) );
OAI211_X2 \myreg/_4429_ ( .A(\myreg/_1929_ ), .B(fanout_net_57 ), .C1(\myreg/_0168_ ), .C2(fanout_net_50 ), .ZN(\myreg/_1930_ ) );
AOI21_X1 \myreg/_4430_ ( .A(fanout_net_57 ), .B1(\myreg/_1358_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1931_ ) );
OAI21_X1 \myreg/_4431_ ( .A(\myreg/_1931_ ), .B1(\myreg/_0104_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1932_ ) );
AOI21_X1 \myreg/_4432_ ( .A(\myreg/_1642_ ), .B1(\myreg/_1930_ ), .B2(\myreg/_1932_ ), .ZN(\myreg/_1933_ ) );
OR2_X1 \myreg/_4433_ ( .A1(\myreg/_0040_ ), .A2(fanout_net_50 ), .ZN(\myreg/_1934_ ) );
OAI211_X2 \myreg/_4434_ ( .A(\myreg/_1934_ ), .B(fanout_net_57 ), .C1(\myreg/_0072_ ), .C2(\myreg/_1679_ ), .ZN(\myreg/_1935_ ) );
AOI21_X1 \myreg/_4435_ ( .A(fanout_net_57 ), .B1(\myreg/_1352_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1936_ ) );
OAI21_X1 \myreg/_4436_ ( .A(\myreg/_1936_ ), .B1(\myreg/_0456_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1937_ ) );
AOI21_X1 \myreg/_4437_ ( .A(fanout_net_60 ), .B1(\myreg/_1935_ ), .B2(\myreg/_1937_ ), .ZN(\myreg/_1938_ ) );
OR2_X1 \myreg/_4438_ ( .A1(\myreg/_1933_ ), .A2(\myreg/_1938_ ), .ZN(\myreg/_1939_ ) );
MUX2_X1 \myreg/_4439_ ( .A(\myreg/_0328_ ), .B(\myreg/_0360_ ), .S(fanout_net_50 ), .Z(\myreg/_1940_ ) );
MUX2_X1 \myreg/_4440_ ( .A(\myreg/_0392_ ), .B(\myreg/_0424_ ), .S(fanout_net_50 ), .Z(\myreg/_1941_ ) );
MUX2_X1 \myreg/_4441_ ( .A(\myreg/_1940_ ), .B(\myreg/_1941_ ), .S(fanout_net_57 ), .Z(\myreg/_1942_ ) );
MUX2_X1 \myreg/_4442_ ( .A(\myreg/_0008_ ), .B(\myreg/_0232_ ), .S(fanout_net_50 ), .Z(\myreg/_1943_ ) );
MUX2_X1 \myreg/_4443_ ( .A(\myreg/_0264_ ), .B(\myreg/_0296_ ), .S(fanout_net_50 ), .Z(\myreg/_1944_ ) );
MUX2_X1 \myreg/_4444_ ( .A(\myreg/_1943_ ), .B(\myreg/_1944_ ), .S(fanout_net_57 ), .Z(\myreg/_1945_ ) );
MUX2_X1 \myreg/_4445_ ( .A(\myreg/_1942_ ), .B(\myreg/_1945_ ), .S(\myreg/_1895_ ), .Z(\myreg/_1946_ ) );
MUX2_X1 \myreg/_4446_ ( .A(\myreg/_1939_ ), .B(\myreg/_1946_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2388_ ) );
OR2_X1 \myreg/_4447_ ( .A1(\myreg/_1679_ ), .A2(\myreg/_0201_ ), .ZN(\myreg/_1947_ ) );
OAI211_X2 \myreg/_4448_ ( .A(\myreg/_1947_ ), .B(fanout_net_57 ), .C1(\myreg/_0169_ ), .C2(fanout_net_50 ), .ZN(\myreg/_1948_ ) );
AOI21_X1 \myreg/_4449_ ( .A(fanout_net_57 ), .B1(\myreg/_1372_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1949_ ) );
OAI21_X1 \myreg/_4450_ ( .A(\myreg/_1949_ ), .B1(\myreg/_0105_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1950_ ) );
NAND3_X1 \myreg/_4451_ ( .A1(\myreg/_1948_ ), .A2(fanout_net_60 ), .A3(\myreg/_1950_ ), .ZN(\myreg/_1951_ ) );
OR2_X1 \myreg/_4452_ ( .A1(\myreg/_1635_ ), .A2(\myreg/_0073_ ), .ZN(\myreg/_1952_ ) );
OAI211_X2 \myreg/_4453_ ( .A(\myreg/_1952_ ), .B(fanout_net_57 ), .C1(\myreg/_0041_ ), .C2(fanout_net_50 ), .ZN(\myreg/_1953_ ) );
AOI21_X1 \myreg/_4454_ ( .A(fanout_net_57 ), .B1(\myreg/_1378_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1954_ ) );
OAI21_X1 \myreg/_4455_ ( .A(\myreg/_1954_ ), .B1(\myreg/_0457_ ), .B2(fanout_net_50 ), .ZN(\myreg/_1955_ ) );
NAND3_X1 \myreg/_4456_ ( .A1(\myreg/_1953_ ), .A2(\myreg/_1656_ ), .A3(\myreg/_1955_ ), .ZN(\myreg/_1956_ ) );
AND2_X1 \myreg/_4457_ ( .A1(\myreg/_1951_ ), .A2(\myreg/_1956_ ), .ZN(\myreg/_1957_ ) );
MUX2_X1 \myreg/_4458_ ( .A(\myreg/_0329_ ), .B(\myreg/_0361_ ), .S(fanout_net_50 ), .Z(\myreg/_1958_ ) );
MUX2_X1 \myreg/_4459_ ( .A(\myreg/_0393_ ), .B(\myreg/_0425_ ), .S(fanout_net_50 ), .Z(\myreg/_1959_ ) );
MUX2_X1 \myreg/_4460_ ( .A(\myreg/_1958_ ), .B(\myreg/_1959_ ), .S(fanout_net_57 ), .Z(\myreg/_1960_ ) );
MUX2_X1 \myreg/_4461_ ( .A(\myreg/_0009_ ), .B(\myreg/_0233_ ), .S(fanout_net_50 ), .Z(\myreg/_1961_ ) );
MUX2_X1 \myreg/_4462_ ( .A(\myreg/_0265_ ), .B(\myreg/_0297_ ), .S(fanout_net_50 ), .Z(\myreg/_1962_ ) );
MUX2_X1 \myreg/_4463_ ( .A(\myreg/_1961_ ), .B(\myreg/_1962_ ), .S(fanout_net_57 ), .Z(\myreg/_1963_ ) );
MUX2_X1 \myreg/_4464_ ( .A(\myreg/_1960_ ), .B(\myreg/_1963_ ), .S(\myreg/_1895_ ), .Z(\myreg/_1964_ ) );
MUX2_X1 \myreg/_4465_ ( .A(\myreg/_1957_ ), .B(\myreg/_1964_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2389_ ) );
MUX2_X1 \myreg/_4466_ ( .A(\myreg/_0106_ ), .B(\myreg/_0138_ ), .S(fanout_net_50 ), .Z(\myreg/_1965_ ) );
MUX2_X1 \myreg/_4467_ ( .A(\myreg/_0170_ ), .B(\myreg/_0202_ ), .S(fanout_net_50 ), .Z(\myreg/_1966_ ) );
MUX2_X1 \myreg/_4468_ ( .A(\myreg/_1965_ ), .B(\myreg/_1966_ ), .S(fanout_net_57 ), .Z(\myreg/_1967_ ) );
MUX2_X1 \myreg/_4469_ ( .A(\myreg/_0458_ ), .B(\myreg/_0490_ ), .S(fanout_net_50 ), .Z(\myreg/_1968_ ) );
MUX2_X1 \myreg/_4470_ ( .A(\myreg/_0042_ ), .B(\myreg/_0074_ ), .S(fanout_net_51 ), .Z(\myreg/_1969_ ) );
MUX2_X1 \myreg/_4471_ ( .A(\myreg/_1968_ ), .B(\myreg/_1969_ ), .S(fanout_net_57 ), .Z(\myreg/_1970_ ) );
MUX2_X1 \myreg/_4472_ ( .A(\myreg/_1967_ ), .B(\myreg/_1970_ ), .S(\myreg/_1660_ ), .Z(\myreg/_1971_ ) );
MUX2_X1 \myreg/_4473_ ( .A(\myreg/_0010_ ), .B(\myreg/_0266_ ), .S(fanout_net_57 ), .Z(\myreg/_1972_ ) );
MUX2_X1 \myreg/_4474_ ( .A(\myreg/_0234_ ), .B(\myreg/_0298_ ), .S(fanout_net_57 ), .Z(\myreg/_1973_ ) );
MUX2_X1 \myreg/_4475_ ( .A(\myreg/_1972_ ), .B(\myreg/_1973_ ), .S(fanout_net_51 ), .Z(\myreg/_1974_ ) );
MUX2_X1 \myreg/_4476_ ( .A(\myreg/_0330_ ), .B(\myreg/_0394_ ), .S(fanout_net_57 ), .Z(\myreg/_1975_ ) );
MUX2_X1 \myreg/_4477_ ( .A(\myreg/_0362_ ), .B(\myreg/_0426_ ), .S(fanout_net_57 ), .Z(\myreg/_1976_ ) );
MUX2_X1 \myreg/_4478_ ( .A(\myreg/_1975_ ), .B(\myreg/_1976_ ), .S(fanout_net_51 ), .Z(\myreg/_1977_ ) );
MUX2_X1 \myreg/_4479_ ( .A(\myreg/_1974_ ), .B(\myreg/_1977_ ), .S(fanout_net_60 ), .Z(\myreg/_1978_ ) );
MUX2_X1 \myreg/_4480_ ( .A(\myreg/_1971_ ), .B(\myreg/_1978_ ), .S(\myreg/_1831_ ), .Z(\myreg/_2390_ ) );
MUX2_X1 \myreg/_4481_ ( .A(\myreg/_0108_ ), .B(\myreg/_0140_ ), .S(fanout_net_51 ), .Z(\myreg/_1979_ ) );
MUX2_X1 \myreg/_4482_ ( .A(\myreg/_0172_ ), .B(\myreg/_0204_ ), .S(fanout_net_51 ), .Z(\myreg/_1980_ ) );
MUX2_X1 \myreg/_4483_ ( .A(\myreg/_1979_ ), .B(\myreg/_1980_ ), .S(fanout_net_57 ), .Z(\myreg/_1981_ ) );
MUX2_X1 \myreg/_4484_ ( .A(\myreg/_0460_ ), .B(\myreg/_0492_ ), .S(fanout_net_51 ), .Z(\myreg/_1982_ ) );
MUX2_X1 \myreg/_4485_ ( .A(\myreg/_0044_ ), .B(\myreg/_0076_ ), .S(fanout_net_51 ), .Z(\myreg/_1983_ ) );
MUX2_X1 \myreg/_4486_ ( .A(\myreg/_1982_ ), .B(\myreg/_1983_ ), .S(fanout_net_57 ), .Z(\myreg/_1984_ ) );
MUX2_X1 \myreg/_4487_ ( .A(\myreg/_1981_ ), .B(\myreg/_1984_ ), .S(\myreg/_1660_ ), .Z(\myreg/_1985_ ) );
MUX2_X1 \myreg/_4488_ ( .A(\myreg/_0012_ ), .B(\myreg/_0268_ ), .S(fanout_net_57 ), .Z(\myreg/_1986_ ) );
MUX2_X1 \myreg/_4489_ ( .A(\myreg/_0236_ ), .B(\myreg/_0300_ ), .S(fanout_net_57 ), .Z(\myreg/_1987_ ) );
MUX2_X1 \myreg/_4490_ ( .A(\myreg/_1986_ ), .B(\myreg/_1987_ ), .S(fanout_net_51 ), .Z(\myreg/_1988_ ) );
MUX2_X1 \myreg/_4491_ ( .A(\myreg/_0332_ ), .B(\myreg/_0396_ ), .S(fanout_net_57 ), .Z(\myreg/_1989_ ) );
MUX2_X1 \myreg/_4492_ ( .A(\myreg/_0364_ ), .B(\myreg/_0428_ ), .S(fanout_net_57 ), .Z(\myreg/_1990_ ) );
MUX2_X1 \myreg/_4493_ ( .A(\myreg/_1989_ ), .B(\myreg/_1990_ ), .S(fanout_net_51 ), .Z(\myreg/_1991_ ) );
MUX2_X1 \myreg/_4494_ ( .A(\myreg/_1988_ ), .B(\myreg/_1991_ ), .S(fanout_net_60 ), .Z(\myreg/_1992_ ) );
BUF_X4 \myreg/_4495_ ( .A(\myreg/_1658_ ), .Z(\myreg/_1993_ ) );
MUX2_X1 \myreg/_4496_ ( .A(\myreg/_1985_ ), .B(\myreg/_1992_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2392_ ) );
MUX2_X1 \myreg/_4497_ ( .A(\myreg/_0109_ ), .B(\myreg/_0141_ ), .S(fanout_net_51 ), .Z(\myreg/_1994_ ) );
MUX2_X1 \myreg/_4498_ ( .A(\myreg/_0173_ ), .B(\myreg/_0205_ ), .S(fanout_net_51 ), .Z(\myreg/_1995_ ) );
MUX2_X1 \myreg/_4499_ ( .A(\myreg/_1994_ ), .B(\myreg/_1995_ ), .S(fanout_net_57 ), .Z(\myreg/_1996_ ) );
MUX2_X1 \myreg/_4500_ ( .A(\myreg/_0461_ ), .B(\myreg/_0493_ ), .S(fanout_net_51 ), .Z(\myreg/_1997_ ) );
MUX2_X1 \myreg/_4501_ ( .A(\myreg/_0045_ ), .B(\myreg/_0077_ ), .S(fanout_net_51 ), .Z(\myreg/_1998_ ) );
MUX2_X1 \myreg/_4502_ ( .A(\myreg/_1997_ ), .B(\myreg/_1998_ ), .S(fanout_net_57 ), .Z(\myreg/_1999_ ) );
MUX2_X1 \myreg/_4503_ ( .A(\myreg/_1996_ ), .B(\myreg/_1999_ ), .S(\myreg/_1660_ ), .Z(\myreg/_2000_ ) );
MUX2_X1 \myreg/_4504_ ( .A(\myreg/_0013_ ), .B(\myreg/_0269_ ), .S(fanout_net_57 ), .Z(\myreg/_2001_ ) );
MUX2_X1 \myreg/_4505_ ( .A(\myreg/_0237_ ), .B(\myreg/_0301_ ), .S(fanout_net_57 ), .Z(\myreg/_2002_ ) );
MUX2_X1 \myreg/_4506_ ( .A(\myreg/_2001_ ), .B(\myreg/_2002_ ), .S(fanout_net_51 ), .Z(\myreg/_2003_ ) );
MUX2_X1 \myreg/_4507_ ( .A(\myreg/_0333_ ), .B(\myreg/_0397_ ), .S(fanout_net_58 ), .Z(\myreg/_2004_ ) );
MUX2_X1 \myreg/_4508_ ( .A(\myreg/_0365_ ), .B(\myreg/_0429_ ), .S(fanout_net_58 ), .Z(\myreg/_2005_ ) );
MUX2_X1 \myreg/_4509_ ( .A(\myreg/_2004_ ), .B(\myreg/_2005_ ), .S(fanout_net_51 ), .Z(\myreg/_2006_ ) );
MUX2_X1 \myreg/_4510_ ( .A(\myreg/_2003_ ), .B(\myreg/_2006_ ), .S(fanout_net_60 ), .Z(\myreg/_2007_ ) );
MUX2_X1 \myreg/_4511_ ( .A(\myreg/_2000_ ), .B(\myreg/_2007_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2393_ ) );
OR2_X1 \myreg/_4512_ ( .A1(\myreg/_0174_ ), .A2(fanout_net_51 ), .ZN(\myreg/_2008_ ) );
OAI211_X2 \myreg/_4513_ ( .A(\myreg/_2008_ ), .B(fanout_net_58 ), .C1(\myreg/_0206_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_2009_ ) );
AOI21_X1 \myreg/_4514_ ( .A(fanout_net_58 ), .B1(\myreg/_1460_ ), .B2(fanout_net_51 ), .ZN(\myreg/_2010_ ) );
OAI21_X1 \myreg/_4515_ ( .A(\myreg/_2010_ ), .B1(\myreg/_0110_ ), .B2(fanout_net_51 ), .ZN(\myreg/_2011_ ) );
NAND3_X1 \myreg/_4516_ ( .A1(\myreg/_2009_ ), .A2(\myreg/_2011_ ), .A3(fanout_net_60 ), .ZN(\myreg/_2012_ ) );
OR2_X1 \myreg/_4517_ ( .A1(\myreg/_0046_ ), .A2(fanout_net_51 ), .ZN(\myreg/_2013_ ) );
OAI211_X2 \myreg/_4518_ ( .A(\myreg/_2013_ ), .B(fanout_net_58 ), .C1(\myreg/_0078_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_2014_ ) );
AOI21_X1 \myreg/_4519_ ( .A(fanout_net_58 ), .B1(\myreg/_1454_ ), .B2(fanout_net_51 ), .ZN(\myreg/_2015_ ) );
OAI21_X1 \myreg/_4520_ ( .A(\myreg/_2015_ ), .B1(\myreg/_0462_ ), .B2(fanout_net_51 ), .ZN(\myreg/_2016_ ) );
NAND3_X1 \myreg/_4521_ ( .A1(\myreg/_2014_ ), .A2(\myreg/_2016_ ), .A3(\myreg/_1656_ ), .ZN(\myreg/_2017_ ) );
AND2_X1 \myreg/_4522_ ( .A1(\myreg/_2012_ ), .A2(\myreg/_2017_ ), .ZN(\myreg/_2018_ ) );
MUX2_X1 \myreg/_4523_ ( .A(\myreg/_0334_ ), .B(\myreg/_0366_ ), .S(fanout_net_51 ), .Z(\myreg/_2019_ ) );
MUX2_X1 \myreg/_4524_ ( .A(\myreg/_0398_ ), .B(\myreg/_0430_ ), .S(fanout_net_51 ), .Z(\myreg/_2020_ ) );
MUX2_X1 \myreg/_4525_ ( .A(\myreg/_2019_ ), .B(\myreg/_2020_ ), .S(fanout_net_58 ), .Z(\myreg/_2021_ ) );
MUX2_X1 \myreg/_4526_ ( .A(\myreg/_0014_ ), .B(\myreg/_0238_ ), .S(fanout_net_51 ), .Z(\myreg/_2022_ ) );
MUX2_X1 \myreg/_4527_ ( .A(\myreg/_0270_ ), .B(\myreg/_0302_ ), .S(fanout_net_51 ), .Z(\myreg/_2023_ ) );
MUX2_X1 \myreg/_4528_ ( .A(\myreg/_2022_ ), .B(\myreg/_2023_ ), .S(fanout_net_58 ), .Z(\myreg/_2024_ ) );
MUX2_X1 \myreg/_4529_ ( .A(\myreg/_2021_ ), .B(\myreg/_2024_ ), .S(\myreg/_1895_ ), .Z(\myreg/_2025_ ) );
MUX2_X1 \myreg/_4530_ ( .A(\myreg/_2018_ ), .B(\myreg/_2025_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2394_ ) );
MUX2_X1 \myreg/_4531_ ( .A(\myreg/_0463_ ), .B(\myreg/_0495_ ), .S(fanout_net_51 ), .Z(\myreg/_2026_ ) );
MUX2_X1 \myreg/_4532_ ( .A(\myreg/_0047_ ), .B(\myreg/_0079_ ), .S(fanout_net_51 ), .Z(\myreg/_2027_ ) );
MUX2_X1 \myreg/_4533_ ( .A(\myreg/_2026_ ), .B(\myreg/_2027_ ), .S(fanout_net_58 ), .Z(\myreg/_2028_ ) );
MUX2_X1 \myreg/_4534_ ( .A(\myreg/_0111_ ), .B(\myreg/_0143_ ), .S(fanout_net_51 ), .Z(\myreg/_2029_ ) );
MUX2_X1 \myreg/_4535_ ( .A(\myreg/_0175_ ), .B(\myreg/_0207_ ), .S(fanout_net_51 ), .Z(\myreg/_2030_ ) );
MUX2_X1 \myreg/_4536_ ( .A(\myreg/_2029_ ), .B(\myreg/_2030_ ), .S(fanout_net_58 ), .Z(\myreg/_2031_ ) );
MUX2_X1 \myreg/_4537_ ( .A(\myreg/_2028_ ), .B(\myreg/_2031_ ), .S(fanout_net_60 ), .Z(\myreg/_2032_ ) );
MUX2_X1 \myreg/_4538_ ( .A(\myreg/_0335_ ), .B(\myreg/_0367_ ), .S(fanout_net_51 ), .Z(\myreg/_2033_ ) );
MUX2_X1 \myreg/_4539_ ( .A(\myreg/_0399_ ), .B(\myreg/_0431_ ), .S(fanout_net_52 ), .Z(\myreg/_2034_ ) );
MUX2_X1 \myreg/_4540_ ( .A(\myreg/_2033_ ), .B(\myreg/_2034_ ), .S(fanout_net_58 ), .Z(\myreg/_2035_ ) );
MUX2_X1 \myreg/_4541_ ( .A(\myreg/_0015_ ), .B(\myreg/_0239_ ), .S(fanout_net_52 ), .Z(\myreg/_2036_ ) );
MUX2_X1 \myreg/_4542_ ( .A(\myreg/_0271_ ), .B(\myreg/_0303_ ), .S(fanout_net_52 ), .Z(\myreg/_2037_ ) );
MUX2_X1 \myreg/_4543_ ( .A(\myreg/_2036_ ), .B(\myreg/_2037_ ), .S(fanout_net_58 ), .Z(\myreg/_2038_ ) );
MUX2_X1 \myreg/_4544_ ( .A(\myreg/_2035_ ), .B(\myreg/_2038_ ), .S(\myreg/_1895_ ), .Z(\myreg/_2039_ ) );
MUX2_X1 \myreg/_4545_ ( .A(\myreg/_2032_ ), .B(\myreg/_2039_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2395_ ) );
MUX2_X1 \myreg/_4546_ ( .A(\myreg/_0112_ ), .B(\myreg/_0144_ ), .S(fanout_net_52 ), .Z(\myreg/_2040_ ) );
MUX2_X1 \myreg/_4547_ ( .A(\myreg/_0176_ ), .B(\myreg/_0208_ ), .S(fanout_net_52 ), .Z(\myreg/_2041_ ) );
MUX2_X1 \myreg/_4548_ ( .A(\myreg/_2040_ ), .B(\myreg/_2041_ ), .S(fanout_net_58 ), .Z(\myreg/_2042_ ) );
MUX2_X1 \myreg/_4549_ ( .A(\myreg/_0464_ ), .B(\myreg/_0496_ ), .S(fanout_net_52 ), .Z(\myreg/_2043_ ) );
MUX2_X1 \myreg/_4550_ ( .A(\myreg/_0048_ ), .B(\myreg/_0080_ ), .S(fanout_net_52 ), .Z(\myreg/_2044_ ) );
MUX2_X1 \myreg/_4551_ ( .A(\myreg/_2043_ ), .B(\myreg/_2044_ ), .S(fanout_net_58 ), .Z(\myreg/_2045_ ) );
MUX2_X1 \myreg/_4552_ ( .A(\myreg/_2042_ ), .B(\myreg/_2045_ ), .S(\myreg/_1660_ ), .Z(\myreg/_2046_ ) );
MUX2_X1 \myreg/_4553_ ( .A(\myreg/_0016_ ), .B(\myreg/_0272_ ), .S(fanout_net_58 ), .Z(\myreg/_2047_ ) );
MUX2_X1 \myreg/_4554_ ( .A(\myreg/_0240_ ), .B(\myreg/_0304_ ), .S(fanout_net_58 ), .Z(\myreg/_2048_ ) );
MUX2_X1 \myreg/_4555_ ( .A(\myreg/_2047_ ), .B(\myreg/_2048_ ), .S(fanout_net_52 ), .Z(\myreg/_2049_ ) );
MUX2_X1 \myreg/_4556_ ( .A(\myreg/_0336_ ), .B(\myreg/_0400_ ), .S(fanout_net_58 ), .Z(\myreg/_2050_ ) );
MUX2_X1 \myreg/_4557_ ( .A(\myreg/_0368_ ), .B(\myreg/_0432_ ), .S(fanout_net_58 ), .Z(\myreg/_2051_ ) );
MUX2_X1 \myreg/_4558_ ( .A(\myreg/_2050_ ), .B(\myreg/_2051_ ), .S(fanout_net_52 ), .Z(\myreg/_2052_ ) );
MUX2_X1 \myreg/_4559_ ( .A(\myreg/_2049_ ), .B(\myreg/_2052_ ), .S(fanout_net_60 ), .Z(\myreg/_2053_ ) );
MUX2_X1 \myreg/_4560_ ( .A(\myreg/_2046_ ), .B(\myreg/_2053_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2396_ ) );
MUX2_X1 \myreg/_4561_ ( .A(\myreg/_0113_ ), .B(\myreg/_0145_ ), .S(fanout_net_52 ), .Z(\myreg/_2054_ ) );
MUX2_X1 \myreg/_4562_ ( .A(\myreg/_0177_ ), .B(\myreg/_0209_ ), .S(fanout_net_52 ), .Z(\myreg/_2055_ ) );
MUX2_X1 \myreg/_4563_ ( .A(\myreg/_2054_ ), .B(\myreg/_2055_ ), .S(fanout_net_58 ), .Z(\myreg/_2056_ ) );
MUX2_X1 \myreg/_4564_ ( .A(\myreg/_0465_ ), .B(\myreg/_0497_ ), .S(fanout_net_52 ), .Z(\myreg/_2057_ ) );
MUX2_X1 \myreg/_4565_ ( .A(\myreg/_0049_ ), .B(\myreg/_0081_ ), .S(fanout_net_52 ), .Z(\myreg/_2058_ ) );
MUX2_X1 \myreg/_4566_ ( .A(\myreg/_2057_ ), .B(\myreg/_2058_ ), .S(fanout_net_58 ), .Z(\myreg/_2059_ ) );
MUX2_X1 \myreg/_4567_ ( .A(\myreg/_2056_ ), .B(\myreg/_2059_ ), .S(\myreg/_1660_ ), .Z(\myreg/_2060_ ) );
MUX2_X1 \myreg/_4568_ ( .A(\myreg/_0017_ ), .B(\myreg/_0273_ ), .S(fanout_net_58 ), .Z(\myreg/_2061_ ) );
MUX2_X1 \myreg/_4569_ ( .A(\myreg/_0241_ ), .B(\myreg/_0305_ ), .S(fanout_net_58 ), .Z(\myreg/_2062_ ) );
MUX2_X1 \myreg/_4570_ ( .A(\myreg/_2061_ ), .B(\myreg/_2062_ ), .S(fanout_net_52 ), .Z(\myreg/_2063_ ) );
MUX2_X1 \myreg/_4571_ ( .A(\myreg/_0337_ ), .B(\myreg/_0401_ ), .S(fanout_net_58 ), .Z(\myreg/_2064_ ) );
MUX2_X1 \myreg/_4572_ ( .A(\myreg/_0369_ ), .B(\myreg/_0433_ ), .S(fanout_net_58 ), .Z(\myreg/_2065_ ) );
MUX2_X1 \myreg/_4573_ ( .A(\myreg/_2064_ ), .B(\myreg/_2065_ ), .S(fanout_net_52 ), .Z(\myreg/_2066_ ) );
MUX2_X1 \myreg/_4574_ ( .A(\myreg/_2063_ ), .B(\myreg/_2066_ ), .S(fanout_net_60 ), .Z(\myreg/_2067_ ) );
MUX2_X1 \myreg/_4575_ ( .A(\myreg/_2060_ ), .B(\myreg/_2067_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2397_ ) );
OR2_X1 \myreg/_4576_ ( .A1(\myreg/_1679_ ), .A2(\myreg/_0082_ ), .ZN(\myreg/_2068_ ) );
OAI211_X2 \myreg/_4577_ ( .A(\myreg/_2068_ ), .B(fanout_net_58 ), .C1(\myreg/_0050_ ), .C2(fanout_net_52 ), .ZN(\myreg/_2069_ ) );
AOI21_X1 \myreg/_4578_ ( .A(fanout_net_58 ), .B1(\myreg/_1534_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2070_ ) );
OAI21_X1 \myreg/_4579_ ( .A(\myreg/_2070_ ), .B1(\myreg/_0466_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2071_ ) );
NAND3_X1 \myreg/_4580_ ( .A1(\myreg/_2069_ ), .A2(\myreg/_1656_ ), .A3(\myreg/_2071_ ), .ZN(\myreg/_2072_ ) );
OR2_X1 \myreg/_4581_ ( .A1(\myreg/_0178_ ), .A2(fanout_net_52 ), .ZN(\myreg/_2073_ ) );
OAI211_X2 \myreg/_4582_ ( .A(\myreg/_2073_ ), .B(fanout_net_58 ), .C1(\myreg/_0210_ ), .C2(\myreg/_1644_ ), .ZN(\myreg/_2074_ ) );
AOI21_X1 \myreg/_4583_ ( .A(fanout_net_58 ), .B1(\myreg/_1528_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2075_ ) );
OAI21_X1 \myreg/_4584_ ( .A(\myreg/_2075_ ), .B1(\myreg/_0114_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2076_ ) );
NAND3_X1 \myreg/_4585_ ( .A1(\myreg/_2074_ ), .A2(\myreg/_2076_ ), .A3(fanout_net_60 ), .ZN(\myreg/_2077_ ) );
AND2_X1 \myreg/_4586_ ( .A1(\myreg/_2072_ ), .A2(\myreg/_2077_ ), .ZN(\myreg/_2078_ ) );
MUX2_X1 \myreg/_4587_ ( .A(\myreg/_0338_ ), .B(\myreg/_0370_ ), .S(fanout_net_52 ), .Z(\myreg/_2079_ ) );
MUX2_X1 \myreg/_4588_ ( .A(\myreg/_0402_ ), .B(\myreg/_0434_ ), .S(fanout_net_52 ), .Z(\myreg/_2080_ ) );
MUX2_X1 \myreg/_4589_ ( .A(\myreg/_2079_ ), .B(\myreg/_2080_ ), .S(fanout_net_58 ), .Z(\myreg/_2081_ ) );
MUX2_X1 \myreg/_4590_ ( .A(\myreg/_0018_ ), .B(\myreg/_0242_ ), .S(fanout_net_52 ), .Z(\myreg/_2082_ ) );
MUX2_X1 \myreg/_4591_ ( .A(\myreg/_0274_ ), .B(\myreg/_0306_ ), .S(fanout_net_52 ), .Z(\myreg/_2083_ ) );
MUX2_X1 \myreg/_4592_ ( .A(\myreg/_2082_ ), .B(\myreg/_2083_ ), .S(fanout_net_58 ), .Z(\myreg/_2084_ ) );
MUX2_X1 \myreg/_4593_ ( .A(\myreg/_2081_ ), .B(\myreg/_2084_ ), .S(\myreg/_1895_ ), .Z(\myreg/_2085_ ) );
MUX2_X1 \myreg/_4594_ ( .A(\myreg/_2078_ ), .B(\myreg/_2085_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2398_ ) );
OR2_X1 \myreg/_4595_ ( .A1(\myreg/_1634_ ), .A2(\myreg/_0083_ ), .ZN(\myreg/_2086_ ) );
OAI211_X2 \myreg/_4596_ ( .A(\myreg/_2086_ ), .B(fanout_net_59 ), .C1(\myreg/_0051_ ), .C2(fanout_net_52 ), .ZN(\myreg/_2087_ ) );
AOI21_X1 \myreg/_4597_ ( .A(fanout_net_59 ), .B1(\myreg/_1548_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2088_ ) );
OAI21_X1 \myreg/_4598_ ( .A(\myreg/_2088_ ), .B1(\myreg/_0467_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2089_ ) );
AOI21_X1 \myreg/_4599_ ( .A(fanout_net_60 ), .B1(\myreg/_2087_ ), .B2(\myreg/_2089_ ), .ZN(\myreg/_2090_ ) );
OR2_X1 \myreg/_4600_ ( .A1(\myreg/_0179_ ), .A2(fanout_net_52 ), .ZN(\myreg/_2091_ ) );
OAI211_X2 \myreg/_4601_ ( .A(\myreg/_2091_ ), .B(fanout_net_59 ), .C1(\myreg/_0211_ ), .C2(\myreg/_1679_ ), .ZN(\myreg/_2092_ ) );
AOI21_X1 \myreg/_4602_ ( .A(fanout_net_59 ), .B1(\myreg/_1554_ ), .B2(fanout_net_52 ), .ZN(\myreg/_2093_ ) );
OAI21_X1 \myreg/_4603_ ( .A(\myreg/_2093_ ), .B1(\myreg/_0115_ ), .B2(fanout_net_53 ), .ZN(\myreg/_2094_ ) );
AOI21_X1 \myreg/_4604_ ( .A(\myreg/_1642_ ), .B1(\myreg/_2092_ ), .B2(\myreg/_2094_ ), .ZN(\myreg/_2095_ ) );
OR2_X1 \myreg/_4605_ ( .A1(\myreg/_2090_ ), .A2(\myreg/_2095_ ), .ZN(\myreg/_2096_ ) );
MUX2_X1 \myreg/_4606_ ( .A(\myreg/_0339_ ), .B(\myreg/_0371_ ), .S(fanout_net_53 ), .Z(\myreg/_2097_ ) );
MUX2_X1 \myreg/_4607_ ( .A(\myreg/_0403_ ), .B(\myreg/_0435_ ), .S(fanout_net_53 ), .Z(\myreg/_2098_ ) );
MUX2_X1 \myreg/_4608_ ( .A(\myreg/_2097_ ), .B(\myreg/_2098_ ), .S(fanout_net_59 ), .Z(\myreg/_2099_ ) );
MUX2_X1 \myreg/_4609_ ( .A(\myreg/_0019_ ), .B(\myreg/_0243_ ), .S(fanout_net_53 ), .Z(\myreg/_2100_ ) );
MUX2_X1 \myreg/_4610_ ( .A(\myreg/_0275_ ), .B(\myreg/_0307_ ), .S(fanout_net_53 ), .Z(\myreg/_2101_ ) );
MUX2_X1 \myreg/_4611_ ( .A(\myreg/_2100_ ), .B(\myreg/_2101_ ), .S(fanout_net_59 ), .Z(\myreg/_2102_ ) );
MUX2_X1 \myreg/_4612_ ( .A(\myreg/_2099_ ), .B(\myreg/_2102_ ), .S(\myreg/_1895_ ), .Z(\myreg/_2103_ ) );
MUX2_X1 \myreg/_4613_ ( .A(\myreg/_2096_ ), .B(\myreg/_2103_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2399_ ) );
MUX2_X1 \myreg/_4614_ ( .A(\myreg/_0116_ ), .B(\myreg/_0148_ ), .S(fanout_net_53 ), .Z(\myreg/_2104_ ) );
MUX2_X1 \myreg/_4615_ ( .A(\myreg/_0180_ ), .B(\myreg/_0212_ ), .S(fanout_net_53 ), .Z(\myreg/_2105_ ) );
MUX2_X1 \myreg/_4616_ ( .A(\myreg/_2104_ ), .B(\myreg/_2105_ ), .S(fanout_net_59 ), .Z(\myreg/_2106_ ) );
MUX2_X1 \myreg/_4617_ ( .A(\myreg/_0468_ ), .B(\myreg/_0500_ ), .S(fanout_net_53 ), .Z(\myreg/_2107_ ) );
MUX2_X1 \myreg/_4618_ ( .A(\myreg/_0052_ ), .B(\myreg/_0084_ ), .S(fanout_net_53 ), .Z(\myreg/_2108_ ) );
MUX2_X1 \myreg/_4619_ ( .A(\myreg/_2107_ ), .B(\myreg/_2108_ ), .S(fanout_net_59 ), .Z(\myreg/_2109_ ) );
MUX2_X1 \myreg/_4620_ ( .A(\myreg/_2106_ ), .B(\myreg/_2109_ ), .S(\myreg/_1660_ ), .Z(\myreg/_2110_ ) );
MUX2_X1 \myreg/_4621_ ( .A(\myreg/_0020_ ), .B(\myreg/_0276_ ), .S(fanout_net_59 ), .Z(\myreg/_2111_ ) );
MUX2_X1 \myreg/_4622_ ( .A(\myreg/_0244_ ), .B(\myreg/_0308_ ), .S(fanout_net_59 ), .Z(\myreg/_2112_ ) );
MUX2_X1 \myreg/_4623_ ( .A(\myreg/_2111_ ), .B(\myreg/_2112_ ), .S(fanout_net_53 ), .Z(\myreg/_2113_ ) );
MUX2_X1 \myreg/_4624_ ( .A(\myreg/_0340_ ), .B(\myreg/_0404_ ), .S(fanout_net_59 ), .Z(\myreg/_2114_ ) );
MUX2_X1 \myreg/_4625_ ( .A(\myreg/_0372_ ), .B(\myreg/_0436_ ), .S(fanout_net_59 ), .Z(\myreg/_2115_ ) );
MUX2_X1 \myreg/_4626_ ( .A(\myreg/_2114_ ), .B(\myreg/_2115_ ), .S(fanout_net_53 ), .Z(\myreg/_2116_ ) );
MUX2_X1 \myreg/_4627_ ( .A(\myreg/_2113_ ), .B(\myreg/_2116_ ), .S(fanout_net_60 ), .Z(\myreg/_2117_ ) );
MUX2_X1 \myreg/_4628_ ( .A(\myreg/_2110_ ), .B(\myreg/_2117_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2400_ ) );
MUX2_X1 \myreg/_4629_ ( .A(\myreg/_0117_ ), .B(\myreg/_0149_ ), .S(fanout_net_53 ), .Z(\myreg/_2118_ ) );
MUX2_X1 \myreg/_4630_ ( .A(\myreg/_0181_ ), .B(\myreg/_0213_ ), .S(fanout_net_53 ), .Z(\myreg/_2119_ ) );
MUX2_X1 \myreg/_4631_ ( .A(\myreg/_2118_ ), .B(\myreg/_2119_ ), .S(fanout_net_59 ), .Z(\myreg/_2120_ ) );
MUX2_X1 \myreg/_4632_ ( .A(\myreg/_0469_ ), .B(\myreg/_0501_ ), .S(fanout_net_53 ), .Z(\myreg/_2121_ ) );
MUX2_X1 \myreg/_4633_ ( .A(\myreg/_0053_ ), .B(\myreg/_0085_ ), .S(fanout_net_53 ), .Z(\myreg/_2122_ ) );
MUX2_X1 \myreg/_4634_ ( .A(\myreg/_2121_ ), .B(\myreg/_2122_ ), .S(fanout_net_59 ), .Z(\myreg/_2123_ ) );
MUX2_X1 \myreg/_4635_ ( .A(\myreg/_2120_ ), .B(\myreg/_2123_ ), .S(\myreg/_1660_ ), .Z(\myreg/_2124_ ) );
MUX2_X1 \myreg/_4636_ ( .A(\myreg/_0021_ ), .B(\myreg/_0277_ ), .S(fanout_net_59 ), .Z(\myreg/_2125_ ) );
MUX2_X1 \myreg/_4637_ ( .A(\myreg/_0245_ ), .B(\myreg/_0309_ ), .S(fanout_net_59 ), .Z(\myreg/_2126_ ) );
MUX2_X1 \myreg/_4638_ ( .A(\myreg/_2125_ ), .B(\myreg/_2126_ ), .S(fanout_net_53 ), .Z(\myreg/_2127_ ) );
MUX2_X1 \myreg/_4639_ ( .A(\myreg/_0341_ ), .B(\myreg/_0405_ ), .S(fanout_net_59 ), .Z(\myreg/_2128_ ) );
MUX2_X1 \myreg/_4640_ ( .A(\myreg/_0373_ ), .B(\myreg/_0437_ ), .S(fanout_net_59 ), .Z(\myreg/_2129_ ) );
MUX2_X1 \myreg/_4641_ ( .A(\myreg/_2128_ ), .B(\myreg/_2129_ ), .S(fanout_net_53 ), .Z(\myreg/_2130_ ) );
MUX2_X1 \myreg/_4642_ ( .A(\myreg/_2127_ ), .B(\myreg/_2130_ ), .S(\myreg/_2346_ ), .Z(\myreg/_2131_ ) );
MUX2_X1 \myreg/_4643_ ( .A(\myreg/_2124_ ), .B(\myreg/_2131_ ), .S(\myreg/_1993_ ), .Z(\myreg/_2401_ ) );
MUX2_X1 \myreg/_4644_ ( .A(\myreg/_0119_ ), .B(\myreg/_0151_ ), .S(fanout_net_53 ), .Z(\myreg/_2132_ ) );
MUX2_X1 \myreg/_4645_ ( .A(\myreg/_0183_ ), .B(\myreg/_0215_ ), .S(fanout_net_53 ), .Z(\myreg/_2133_ ) );
MUX2_X1 \myreg/_4646_ ( .A(\myreg/_2132_ ), .B(\myreg/_2133_ ), .S(fanout_net_59 ), .Z(\myreg/_2134_ ) );
MUX2_X1 \myreg/_4647_ ( .A(\myreg/_0471_ ), .B(\myreg/_0503_ ), .S(fanout_net_53 ), .Z(\myreg/_2135_ ) );
MUX2_X1 \myreg/_4648_ ( .A(\myreg/_0055_ ), .B(\myreg/_0087_ ), .S(fanout_net_53 ), .Z(\myreg/_2136_ ) );
MUX2_X1 \myreg/_4649_ ( .A(\myreg/_2135_ ), .B(\myreg/_2136_ ), .S(fanout_net_59 ), .Z(\myreg/_2137_ ) );
MUX2_X1 \myreg/_4650_ ( .A(\myreg/_2134_ ), .B(\myreg/_2137_ ), .S(\myreg/_1660_ ), .Z(\myreg/_2138_ ) );
MUX2_X1 \myreg/_4651_ ( .A(\myreg/_0023_ ), .B(\myreg/_0279_ ), .S(fanout_net_59 ), .Z(\myreg/_2139_ ) );
MUX2_X1 \myreg/_4652_ ( .A(\myreg/_0247_ ), .B(\myreg/_0311_ ), .S(fanout_net_59 ), .Z(\myreg/_2140_ ) );
MUX2_X1 \myreg/_4653_ ( .A(\myreg/_2139_ ), .B(\myreg/_2140_ ), .S(fanout_net_53 ), .Z(\myreg/_2141_ ) );
MUX2_X1 \myreg/_4654_ ( .A(\myreg/_0343_ ), .B(\myreg/_0407_ ), .S(fanout_net_59 ), .Z(\myreg/_2142_ ) );
MUX2_X1 \myreg/_4655_ ( .A(\myreg/_0375_ ), .B(\myreg/_0439_ ), .S(fanout_net_59 ), .Z(\myreg/_2143_ ) );
MUX2_X1 \myreg/_4656_ ( .A(\myreg/_2142_ ), .B(\myreg/_2143_ ), .S(fanout_net_53 ), .Z(\myreg/_2144_ ) );
MUX2_X1 \myreg/_4657_ ( .A(\myreg/_2141_ ), .B(\myreg/_2144_ ), .S(\myreg/_2346_ ), .Z(\myreg/_2145_ ) );
MUX2_X1 \myreg/_4658_ ( .A(\myreg/_2138_ ), .B(\myreg/_2145_ ), .S(\myreg/_1658_ ), .Z(\myreg/_2403_ ) );
MUX2_X1 \myreg/_4659_ ( .A(\myreg/_0472_ ), .B(\myreg/_0504_ ), .S(fanout_net_53 ), .Z(\myreg/_2146_ ) );
MUX2_X1 \myreg/_4660_ ( .A(\myreg/_0056_ ), .B(\myreg/_0088_ ), .S(fanout_net_53 ), .Z(\myreg/_2147_ ) );
MUX2_X1 \myreg/_4661_ ( .A(\myreg/_2146_ ), .B(\myreg/_2147_ ), .S(fanout_net_59 ), .Z(\myreg/_2148_ ) );
MUX2_X1 \myreg/_4662_ ( .A(\myreg/_0120_ ), .B(\myreg/_0152_ ), .S(fanout_net_53 ), .Z(\myreg/_2149_ ) );
MUX2_X1 \myreg/_4663_ ( .A(\myreg/_0184_ ), .B(\myreg/_0216_ ), .S(fanout_net_53 ), .Z(\myreg/_2150_ ) );
MUX2_X1 \myreg/_4664_ ( .A(\myreg/_2149_ ), .B(\myreg/_2150_ ), .S(fanout_net_59 ), .Z(\myreg/_2151_ ) );
MUX2_X1 \myreg/_4665_ ( .A(\myreg/_2148_ ), .B(\myreg/_2151_ ), .S(\myreg/_2346_ ), .Z(\myreg/_2152_ ) );
MUX2_X1 \myreg/_4666_ ( .A(\myreg/_0344_ ), .B(\myreg/_0376_ ), .S(fanout_net_53 ), .Z(\myreg/_2153_ ) );
MUX2_X1 \myreg/_4667_ ( .A(\myreg/_0408_ ), .B(\myreg/_0440_ ), .S(fanout_net_53 ), .Z(\myreg/_2154_ ) );
MUX2_X1 \myreg/_4668_ ( .A(\myreg/_2153_ ), .B(\myreg/_2154_ ), .S(fanout_net_59 ), .Z(\myreg/_2155_ ) );
MUX2_X1 \myreg/_4669_ ( .A(\myreg/_0024_ ), .B(\myreg/_0248_ ), .S(fanout_net_53 ), .Z(\myreg/_2156_ ) );
MUX2_X1 \myreg/_4670_ ( .A(\myreg/_0280_ ), .B(\myreg/_0312_ ), .S(\myreg/_2344_ ), .Z(\myreg/_2157_ ) );
MUX2_X1 \myreg/_4671_ ( .A(\myreg/_2156_ ), .B(\myreg/_2157_ ), .S(fanout_net_59 ), .Z(\myreg/_2158_ ) );
MUX2_X1 \myreg/_4672_ ( .A(\myreg/_2155_ ), .B(\myreg/_2158_ ), .S(\myreg/_1895_ ), .Z(\myreg/_2159_ ) );
MUX2_X1 \myreg/_4673_ ( .A(\myreg/_2152_ ), .B(\myreg/_2159_ ), .S(\myreg/_1658_ ), .Z(\myreg/_2404_ ) );
NOR2_X4 \myreg/_4674_ ( .A1(\myreg/_2413_ ), .A2(\myreg/_2416_ ), .ZN(\myreg/_2160_ ) );
INV_X4 \myreg/_4675_ ( .A(\myreg/_2414_ ), .ZN(\myreg/_2161_ ) );
INV_X4 \myreg/_4676_ ( .A(\myreg/_2415_ ), .ZN(\myreg/_2162_ ) );
NAND3_X4 \myreg/_4677_ ( .A1(\myreg/_2160_ ), .A2(\myreg/_2161_ ), .A3(\myreg/_2162_ ), .ZN(\myreg/_2163_ ) );
NAND2_X4 \myreg/_4678_ ( .A1(\myreg/_2163_ ), .A2(\myreg/_2449_ ), .ZN(\myreg/_2164_ ) );
NOR2_X4 \myreg/_4679_ ( .A1(\myreg/_2164_ ), .A2(fanout_net_61 ), .ZN(\myreg/_2165_ ) );
CLKBUF_X2 \myreg/_4680_ ( .A(\myreg/_2165_ ), .Z(\myreg/_2166_ ) );
AND2_X1 \myreg/_4681_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2417_ ), .ZN(\myreg/_2167_ ) );
CLKBUF_X2 \myreg/_4682_ ( .A(\myreg/_2167_ ), .Z(\myreg/_2168_ ) );
AND2_X4 \myreg/_4683_ ( .A1(\myreg/_2165_ ), .A2(\myreg/_2413_ ), .ZN(\myreg/_2169_ ) );
NAND2_X4 \myreg/_4684_ ( .A1(\myreg/_2169_ ), .A2(\myreg/_2414_ ), .ZN(\myreg/_2170_ ) );
AND2_X4 \myreg/_4685_ ( .A1(\myreg/_2165_ ), .A2(\myreg/_2415_ ), .ZN(\myreg/_2171_ ) );
INV_X1 \myreg/_4686_ ( .A(\myreg/_2416_ ), .ZN(\myreg/_2172_ ) );
NAND2_X4 \myreg/_4687_ ( .A1(\myreg/_2171_ ), .A2(\myreg/_2172_ ), .ZN(\myreg/_2173_ ) );
NOR2_X4 \myreg/_4688_ ( .A1(\myreg/_2170_ ), .A2(\myreg/_2173_ ), .ZN(\myreg/_2174_ ) );
BUF_X4 \myreg/_4689_ ( .A(\myreg/_2174_ ), .Z(\myreg/_2175_ ) );
MUX2_X1 \myreg/_4690_ ( .A(\myreg/_0416_ ), .B(\myreg/_2168_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0512_ ) );
AND2_X1 \myreg/_4691_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2428_ ), .ZN(\myreg/_2176_ ) );
CLKBUF_X2 \myreg/_4692_ ( .A(\myreg/_2176_ ), .Z(\myreg/_2177_ ) );
MUX2_X1 \myreg/_4693_ ( .A(\myreg/_0427_ ), .B(\myreg/_2177_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0513_ ) );
AND2_X1 \myreg/_4694_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2439_ ), .ZN(\myreg/_2178_ ) );
CLKBUF_X2 \myreg/_4695_ ( .A(\myreg/_2178_ ), .Z(\myreg/_2179_ ) );
MUX2_X1 \myreg/_4696_ ( .A(\myreg/_0438_ ), .B(\myreg/_2179_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0514_ ) );
AND2_X1 \myreg/_4697_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2442_ ), .ZN(\myreg/_2180_ ) );
CLKBUF_X2 \myreg/_4698_ ( .A(\myreg/_2180_ ), .Z(\myreg/_2181_ ) );
MUX2_X1 \myreg/_4699_ ( .A(\myreg/_0441_ ), .B(\myreg/_2181_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0515_ ) );
AND2_X1 \myreg/_4700_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2443_ ), .ZN(\myreg/_2182_ ) );
CLKBUF_X2 \myreg/_4701_ ( .A(\myreg/_2182_ ), .Z(\myreg/_2183_ ) );
MUX2_X1 \myreg/_4702_ ( .A(\myreg/_0442_ ), .B(\myreg/_2183_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0516_ ) );
AND2_X1 \myreg/_4703_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2444_ ), .ZN(\myreg/_2184_ ) );
CLKBUF_X2 \myreg/_4704_ ( .A(\myreg/_2184_ ), .Z(\myreg/_2185_ ) );
MUX2_X1 \myreg/_4705_ ( .A(\myreg/_0443_ ), .B(\myreg/_2185_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0517_ ) );
AND2_X1 \myreg/_4706_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2445_ ), .ZN(\myreg/_2186_ ) );
CLKBUF_X2 \myreg/_4707_ ( .A(\myreg/_2186_ ), .Z(\myreg/_2187_ ) );
MUX2_X1 \myreg/_4708_ ( .A(\myreg/_0444_ ), .B(\myreg/_2187_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0518_ ) );
AND2_X1 \myreg/_4709_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2446_ ), .ZN(\myreg/_2188_ ) );
CLKBUF_X2 \myreg/_4710_ ( .A(\myreg/_2188_ ), .Z(\myreg/_2189_ ) );
MUX2_X1 \myreg/_4711_ ( .A(\myreg/_0445_ ), .B(\myreg/_2189_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0519_ ) );
AND2_X1 \myreg/_4712_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2447_ ), .ZN(\myreg/_2190_ ) );
CLKBUF_X2 \myreg/_4713_ ( .A(\myreg/_2190_ ), .Z(\myreg/_2191_ ) );
MUX2_X1 \myreg/_4714_ ( .A(\myreg/_0446_ ), .B(\myreg/_2191_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0520_ ) );
AND2_X1 \myreg/_4715_ ( .A1(\myreg/_2166_ ), .A2(\myreg/_2448_ ), .ZN(\myreg/_2192_ ) );
CLKBUF_X2 \myreg/_4716_ ( .A(\myreg/_2192_ ), .Z(\myreg/_2193_ ) );
MUX2_X1 \myreg/_4717_ ( .A(\myreg/_0447_ ), .B(\myreg/_2193_ ), .S(\myreg/_2175_ ), .Z(\myreg/_0521_ ) );
CLKBUF_X2 \myreg/_4718_ ( .A(\myreg/_2165_ ), .Z(\myreg/_2194_ ) );
AND2_X1 \myreg/_4719_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2418_ ), .ZN(\myreg/_2195_ ) );
CLKBUF_X2 \myreg/_4720_ ( .A(\myreg/_2195_ ), .Z(\myreg/_2196_ ) );
BUF_X4 \myreg/_4721_ ( .A(\myreg/_2174_ ), .Z(\myreg/_2197_ ) );
MUX2_X1 \myreg/_4722_ ( .A(\myreg/_0417_ ), .B(\myreg/_2196_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0522_ ) );
AND2_X1 \myreg/_4723_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2419_ ), .ZN(\myreg/_2198_ ) );
CLKBUF_X2 \myreg/_4724_ ( .A(\myreg/_2198_ ), .Z(\myreg/_2199_ ) );
MUX2_X1 \myreg/_4725_ ( .A(\myreg/_0418_ ), .B(\myreg/_2199_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0523_ ) );
AND2_X1 \myreg/_4726_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2420_ ), .ZN(\myreg/_2200_ ) );
CLKBUF_X2 \myreg/_4727_ ( .A(\myreg/_2200_ ), .Z(\myreg/_2201_ ) );
MUX2_X1 \myreg/_4728_ ( .A(\myreg/_0419_ ), .B(\myreg/_2201_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0524_ ) );
AND2_X1 \myreg/_4729_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2421_ ), .ZN(\myreg/_2202_ ) );
CLKBUF_X2 \myreg/_4730_ ( .A(\myreg/_2202_ ), .Z(\myreg/_2203_ ) );
MUX2_X1 \myreg/_4731_ ( .A(\myreg/_0420_ ), .B(\myreg/_2203_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0525_ ) );
AND2_X1 \myreg/_4732_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2422_ ), .ZN(\myreg/_2204_ ) );
CLKBUF_X2 \myreg/_4733_ ( .A(\myreg/_2204_ ), .Z(\myreg/_2205_ ) );
MUX2_X1 \myreg/_4734_ ( .A(\myreg/_0421_ ), .B(\myreg/_2205_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0526_ ) );
AND2_X1 \myreg/_4735_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2423_ ), .ZN(\myreg/_2206_ ) );
CLKBUF_X2 \myreg/_4736_ ( .A(\myreg/_2206_ ), .Z(\myreg/_2207_ ) );
MUX2_X1 \myreg/_4737_ ( .A(\myreg/_0422_ ), .B(\myreg/_2207_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0527_ ) );
AND2_X1 \myreg/_4738_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2424_ ), .ZN(\myreg/_2208_ ) );
CLKBUF_X2 \myreg/_4739_ ( .A(\myreg/_2208_ ), .Z(\myreg/_2209_ ) );
MUX2_X1 \myreg/_4740_ ( .A(\myreg/_0423_ ), .B(\myreg/_2209_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0528_ ) );
AND2_X1 \myreg/_4741_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2425_ ), .ZN(\myreg/_2210_ ) );
CLKBUF_X2 \myreg/_4742_ ( .A(\myreg/_2210_ ), .Z(\myreg/_2211_ ) );
MUX2_X1 \myreg/_4743_ ( .A(\myreg/_0424_ ), .B(\myreg/_2211_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0529_ ) );
AND2_X1 \myreg/_4744_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2426_ ), .ZN(\myreg/_2212_ ) );
CLKBUF_X2 \myreg/_4745_ ( .A(\myreg/_2212_ ), .Z(\myreg/_2213_ ) );
MUX2_X1 \myreg/_4746_ ( .A(\myreg/_0425_ ), .B(\myreg/_2213_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0530_ ) );
AND2_X1 \myreg/_4747_ ( .A1(\myreg/_2194_ ), .A2(\myreg/_2427_ ), .ZN(\myreg/_2214_ ) );
CLKBUF_X2 \myreg/_4748_ ( .A(\myreg/_2214_ ), .Z(\myreg/_2215_ ) );
MUX2_X1 \myreg/_4749_ ( .A(\myreg/_0426_ ), .B(\myreg/_2215_ ), .S(\myreg/_2197_ ), .Z(\myreg/_0531_ ) );
CLKBUF_X2 \myreg/_4750_ ( .A(\myreg/_2165_ ), .Z(\myreg/_2216_ ) );
AND2_X1 \myreg/_4751_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2429_ ), .ZN(\myreg/_2217_ ) );
CLKBUF_X2 \myreg/_4752_ ( .A(\myreg/_2217_ ), .Z(\myreg/_2218_ ) );
BUF_X4 \myreg/_4753_ ( .A(\myreg/_2174_ ), .Z(\myreg/_2219_ ) );
MUX2_X1 \myreg/_4754_ ( .A(\myreg/_0428_ ), .B(\myreg/_2218_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0532_ ) );
AND2_X1 \myreg/_4755_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2430_ ), .ZN(\myreg/_2220_ ) );
CLKBUF_X2 \myreg/_4756_ ( .A(\myreg/_2220_ ), .Z(\myreg/_2221_ ) );
MUX2_X1 \myreg/_4757_ ( .A(\myreg/_0429_ ), .B(\myreg/_2221_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0533_ ) );
AND2_X1 \myreg/_4758_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2431_ ), .ZN(\myreg/_2222_ ) );
CLKBUF_X2 \myreg/_4759_ ( .A(\myreg/_2222_ ), .Z(\myreg/_2223_ ) );
MUX2_X1 \myreg/_4760_ ( .A(\myreg/_0430_ ), .B(\myreg/_2223_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0534_ ) );
AND2_X1 \myreg/_4761_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2432_ ), .ZN(\myreg/_2224_ ) );
CLKBUF_X2 \myreg/_4762_ ( .A(\myreg/_2224_ ), .Z(\myreg/_2225_ ) );
MUX2_X1 \myreg/_4763_ ( .A(\myreg/_0431_ ), .B(\myreg/_2225_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0535_ ) );
AND2_X1 \myreg/_4764_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2433_ ), .ZN(\myreg/_2226_ ) );
CLKBUF_X2 \myreg/_4765_ ( .A(\myreg/_2226_ ), .Z(\myreg/_2227_ ) );
MUX2_X1 \myreg/_4766_ ( .A(\myreg/_0432_ ), .B(\myreg/_2227_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0536_ ) );
AND2_X1 \myreg/_4767_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2434_ ), .ZN(\myreg/_2228_ ) );
CLKBUF_X2 \myreg/_4768_ ( .A(\myreg/_2228_ ), .Z(\myreg/_2229_ ) );
MUX2_X1 \myreg/_4769_ ( .A(\myreg/_0433_ ), .B(\myreg/_2229_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0537_ ) );
AND2_X1 \myreg/_4770_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2435_ ), .ZN(\myreg/_2230_ ) );
CLKBUF_X2 \myreg/_4771_ ( .A(\myreg/_2230_ ), .Z(\myreg/_2231_ ) );
MUX2_X1 \myreg/_4772_ ( .A(\myreg/_0434_ ), .B(\myreg/_2231_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0538_ ) );
AND2_X1 \myreg/_4773_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2436_ ), .ZN(\myreg/_2232_ ) );
CLKBUF_X2 \myreg/_4774_ ( .A(\myreg/_2232_ ), .Z(\myreg/_2233_ ) );
MUX2_X1 \myreg/_4775_ ( .A(\myreg/_0435_ ), .B(\myreg/_2233_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0539_ ) );
AND2_X1 \myreg/_4776_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2437_ ), .ZN(\myreg/_2234_ ) );
CLKBUF_X2 \myreg/_4777_ ( .A(\myreg/_2234_ ), .Z(\myreg/_2235_ ) );
MUX2_X1 \myreg/_4778_ ( .A(\myreg/_0436_ ), .B(\myreg/_2235_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0540_ ) );
AND2_X1 \myreg/_4779_ ( .A1(\myreg/_2216_ ), .A2(\myreg/_2438_ ), .ZN(\myreg/_2236_ ) );
CLKBUF_X2 \myreg/_4780_ ( .A(\myreg/_2236_ ), .Z(\myreg/_2237_ ) );
MUX2_X1 \myreg/_4781_ ( .A(\myreg/_0437_ ), .B(\myreg/_2237_ ), .S(\myreg/_2219_ ), .Z(\myreg/_0541_ ) );
AND2_X1 \myreg/_4782_ ( .A1(\myreg/_2165_ ), .A2(\myreg/_2440_ ), .ZN(\myreg/_2238_ ) );
CLKBUF_X2 \myreg/_4783_ ( .A(\myreg/_2238_ ), .Z(\myreg/_2239_ ) );
MUX2_X1 \myreg/_4784_ ( .A(\myreg/_0439_ ), .B(\myreg/_2239_ ), .S(\myreg/_2174_ ), .Z(\myreg/_0542_ ) );
AND2_X1 \myreg/_4785_ ( .A1(\myreg/_2165_ ), .A2(\myreg/_2441_ ), .ZN(\myreg/_2240_ ) );
CLKBUF_X2 \myreg/_4786_ ( .A(\myreg/_2240_ ), .Z(\myreg/_2241_ ) );
MUX2_X1 \myreg/_4787_ ( .A(\myreg/_0440_ ), .B(\myreg/_2241_ ), .S(\myreg/_2174_ ), .Z(\myreg/_0543_ ) );
AND2_X2 \myreg/_4788_ ( .A1(\myreg/_2165_ ), .A2(\myreg/_2414_ ), .ZN(\myreg/_2242_ ) );
INV_X1 \myreg/_4789_ ( .A(\myreg/_2413_ ), .ZN(\myreg/_2243_ ) );
NAND2_X4 \myreg/_4790_ ( .A1(\myreg/_2242_ ), .A2(\myreg/_2243_ ), .ZN(\myreg/_2244_ ) );
INV_X2 \myreg/_4791_ ( .A(\myreg/_2165_ ), .ZN(\myreg/_2245_ ) );
AOI21_X4 \myreg/_4792_ ( .A(\myreg/_2245_ ), .B1(\myreg/_2172_ ), .B2(\myreg/_2162_ ), .ZN(\myreg/_2246_ ) );
NOR2_X4 \myreg/_4793_ ( .A1(\myreg/_2244_ ), .A2(\myreg/_2246_ ), .ZN(\myreg/_2247_ ) );
BUF_X8 \myreg/_4794_ ( .A(\myreg/_2247_ ), .Z(\myreg/_2248_ ) );
MUX2_X1 \myreg/_4795_ ( .A(\myreg/_0256_ ), .B(\myreg/_2168_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0544_ ) );
MUX2_X1 \myreg/_4796_ ( .A(\myreg/_0267_ ), .B(\myreg/_2177_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0545_ ) );
MUX2_X1 \myreg/_4797_ ( .A(\myreg/_0278_ ), .B(\myreg/_2179_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0546_ ) );
MUX2_X1 \myreg/_4798_ ( .A(\myreg/_0281_ ), .B(\myreg/_2181_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0547_ ) );
MUX2_X1 \myreg/_4799_ ( .A(\myreg/_0282_ ), .B(\myreg/_2183_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0548_ ) );
MUX2_X1 \myreg/_4800_ ( .A(\myreg/_0283_ ), .B(\myreg/_2185_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0549_ ) );
MUX2_X1 \myreg/_4801_ ( .A(\myreg/_0284_ ), .B(\myreg/_2187_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0550_ ) );
MUX2_X1 \myreg/_4802_ ( .A(\myreg/_0285_ ), .B(\myreg/_2189_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0551_ ) );
MUX2_X1 \myreg/_4803_ ( .A(\myreg/_0286_ ), .B(\myreg/_2191_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0552_ ) );
MUX2_X1 \myreg/_4804_ ( .A(\myreg/_0287_ ), .B(\myreg/_2193_ ), .S(\myreg/_2248_ ), .Z(\myreg/_0553_ ) );
BUF_X8 \myreg/_4805_ ( .A(\myreg/_2247_ ), .Z(\myreg/_2249_ ) );
MUX2_X1 \myreg/_4806_ ( .A(\myreg/_0257_ ), .B(\myreg/_2196_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0554_ ) );
MUX2_X1 \myreg/_4807_ ( .A(\myreg/_0258_ ), .B(\myreg/_2199_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0555_ ) );
MUX2_X1 \myreg/_4808_ ( .A(\myreg/_0259_ ), .B(\myreg/_2201_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0556_ ) );
MUX2_X1 \myreg/_4809_ ( .A(\myreg/_0260_ ), .B(\myreg/_2203_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0557_ ) );
MUX2_X1 \myreg/_4810_ ( .A(\myreg/_0261_ ), .B(\myreg/_2205_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0558_ ) );
MUX2_X1 \myreg/_4811_ ( .A(\myreg/_0262_ ), .B(\myreg/_2207_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0559_ ) );
MUX2_X1 \myreg/_4812_ ( .A(\myreg/_0263_ ), .B(\myreg/_2209_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0560_ ) );
MUX2_X1 \myreg/_4813_ ( .A(\myreg/_0264_ ), .B(\myreg/_2211_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0561_ ) );
MUX2_X1 \myreg/_4814_ ( .A(\myreg/_0265_ ), .B(\myreg/_2213_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0562_ ) );
MUX2_X1 \myreg/_4815_ ( .A(\myreg/_0266_ ), .B(\myreg/_2215_ ), .S(\myreg/_2249_ ), .Z(\myreg/_0563_ ) );
BUF_X8 \myreg/_4816_ ( .A(\myreg/_2247_ ), .Z(\myreg/_2250_ ) );
MUX2_X1 \myreg/_4817_ ( .A(\myreg/_0268_ ), .B(\myreg/_2218_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0564_ ) );
MUX2_X1 \myreg/_4818_ ( .A(\myreg/_0269_ ), .B(\myreg/_2221_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0565_ ) );
MUX2_X1 \myreg/_4819_ ( .A(\myreg/_0270_ ), .B(\myreg/_2223_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0566_ ) );
MUX2_X1 \myreg/_4820_ ( .A(\myreg/_0271_ ), .B(\myreg/_2225_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0567_ ) );
MUX2_X1 \myreg/_4821_ ( .A(\myreg/_0272_ ), .B(\myreg/_2227_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0568_ ) );
MUX2_X1 \myreg/_4822_ ( .A(\myreg/_0273_ ), .B(\myreg/_2229_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0569_ ) );
MUX2_X1 \myreg/_4823_ ( .A(\myreg/_0274_ ), .B(\myreg/_2231_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0570_ ) );
MUX2_X1 \myreg/_4824_ ( .A(\myreg/_0275_ ), .B(\myreg/_2233_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0571_ ) );
MUX2_X1 \myreg/_4825_ ( .A(\myreg/_0276_ ), .B(\myreg/_2235_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0572_ ) );
MUX2_X1 \myreg/_4826_ ( .A(\myreg/_0277_ ), .B(\myreg/_2237_ ), .S(\myreg/_2250_ ), .Z(\myreg/_0573_ ) );
MUX2_X1 \myreg/_4827_ ( .A(\myreg/_0279_ ), .B(\myreg/_2239_ ), .S(\myreg/_2247_ ), .Z(\myreg/_0574_ ) );
MUX2_X1 \myreg/_4828_ ( .A(\myreg/_0280_ ), .B(\myreg/_2241_ ), .S(\myreg/_2247_ ), .Z(\myreg/_0575_ ) );
NAND2_X4 \myreg/_4829_ ( .A1(\myreg/_2169_ ), .A2(\myreg/_2161_ ), .ZN(\myreg/_2251_ ) );
NOR2_X4 \myreg/_4830_ ( .A1(\myreg/_2251_ ), .A2(\myreg/_2246_ ), .ZN(\myreg/_2252_ ) );
BUF_X8 \myreg/_4831_ ( .A(\myreg/_2252_ ), .Z(\myreg/_2253_ ) );
MUX2_X1 \myreg/_4832_ ( .A(\myreg/_0224_ ), .B(\myreg/_2168_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0576_ ) );
MUX2_X1 \myreg/_4833_ ( .A(\myreg/_0235_ ), .B(\myreg/_2177_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0577_ ) );
MUX2_X1 \myreg/_4834_ ( .A(\myreg/_0246_ ), .B(\myreg/_2179_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0578_ ) );
MUX2_X1 \myreg/_4835_ ( .A(\myreg/_0249_ ), .B(\myreg/_2181_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0579_ ) );
MUX2_X1 \myreg/_4836_ ( .A(\myreg/_0250_ ), .B(\myreg/_2183_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0580_ ) );
MUX2_X1 \myreg/_4837_ ( .A(\myreg/_0251_ ), .B(\myreg/_2185_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0581_ ) );
MUX2_X1 \myreg/_4838_ ( .A(\myreg/_0252_ ), .B(\myreg/_2187_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0582_ ) );
MUX2_X1 \myreg/_4839_ ( .A(\myreg/_0253_ ), .B(\myreg/_2189_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0583_ ) );
MUX2_X1 \myreg/_4840_ ( .A(\myreg/_0254_ ), .B(\myreg/_2191_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0584_ ) );
MUX2_X1 \myreg/_4841_ ( .A(\myreg/_0255_ ), .B(\myreg/_2193_ ), .S(\myreg/_2253_ ), .Z(\myreg/_0585_ ) );
BUF_X8 \myreg/_4842_ ( .A(\myreg/_2252_ ), .Z(\myreg/_2254_ ) );
MUX2_X1 \myreg/_4843_ ( .A(\myreg/_0225_ ), .B(\myreg/_2196_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0586_ ) );
MUX2_X1 \myreg/_4844_ ( .A(\myreg/_0226_ ), .B(\myreg/_2199_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0587_ ) );
MUX2_X1 \myreg/_4845_ ( .A(\myreg/_0227_ ), .B(\myreg/_2201_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0588_ ) );
MUX2_X1 \myreg/_4846_ ( .A(\myreg/_0228_ ), .B(\myreg/_2203_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0589_ ) );
MUX2_X1 \myreg/_4847_ ( .A(\myreg/_0229_ ), .B(\myreg/_2205_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0590_ ) );
MUX2_X1 \myreg/_4848_ ( .A(\myreg/_0230_ ), .B(\myreg/_2207_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0591_ ) );
MUX2_X1 \myreg/_4849_ ( .A(\myreg/_0231_ ), .B(\myreg/_2209_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0592_ ) );
MUX2_X1 \myreg/_4850_ ( .A(\myreg/_0232_ ), .B(\myreg/_2211_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0593_ ) );
MUX2_X1 \myreg/_4851_ ( .A(\myreg/_0233_ ), .B(\myreg/_2213_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0594_ ) );
MUX2_X1 \myreg/_4852_ ( .A(\myreg/_0234_ ), .B(\myreg/_2215_ ), .S(\myreg/_2254_ ), .Z(\myreg/_0595_ ) );
BUF_X8 \myreg/_4853_ ( .A(\myreg/_2252_ ), .Z(\myreg/_2255_ ) );
MUX2_X1 \myreg/_4854_ ( .A(\myreg/_0236_ ), .B(\myreg/_2218_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0596_ ) );
MUX2_X1 \myreg/_4855_ ( .A(\myreg/_0237_ ), .B(\myreg/_2221_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0597_ ) );
MUX2_X1 \myreg/_4856_ ( .A(\myreg/_0238_ ), .B(\myreg/_2223_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0598_ ) );
MUX2_X1 \myreg/_4857_ ( .A(\myreg/_0239_ ), .B(\myreg/_2225_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0599_ ) );
MUX2_X1 \myreg/_4858_ ( .A(\myreg/_0240_ ), .B(\myreg/_2227_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0600_ ) );
MUX2_X1 \myreg/_4859_ ( .A(\myreg/_0241_ ), .B(\myreg/_2229_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0601_ ) );
MUX2_X1 \myreg/_4860_ ( .A(\myreg/_0242_ ), .B(\myreg/_2231_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0602_ ) );
MUX2_X1 \myreg/_4861_ ( .A(\myreg/_0243_ ), .B(\myreg/_2233_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0603_ ) );
MUX2_X1 \myreg/_4862_ ( .A(\myreg/_0244_ ), .B(\myreg/_2235_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0604_ ) );
MUX2_X1 \myreg/_4863_ ( .A(\myreg/_0245_ ), .B(\myreg/_2237_ ), .S(\myreg/_2255_ ), .Z(\myreg/_0605_ ) );
MUX2_X1 \myreg/_4864_ ( .A(\myreg/_0247_ ), .B(\myreg/_2239_ ), .S(\myreg/_2252_ ), .Z(\myreg/_0606_ ) );
MUX2_X1 \myreg/_4865_ ( .A(\myreg/_0248_ ), .B(\myreg/_2241_ ), .S(\myreg/_2252_ ), .Z(\myreg/_0607_ ) );
AOI21_X4 \myreg/_4866_ ( .A(\myreg/_2245_ ), .B1(\myreg/_2161_ ), .B2(\myreg/_2243_ ), .ZN(\myreg/_2256_ ) );
NOR2_X4 \myreg/_4867_ ( .A1(\myreg/_2173_ ), .A2(\myreg/_2256_ ), .ZN(\myreg/_2257_ ) );
BUF_X8 \myreg/_4868_ ( .A(\myreg/_2257_ ), .Z(\myreg/_2258_ ) );
MUX2_X1 \myreg/_4869_ ( .A(\myreg/_0320_ ), .B(\myreg/_2168_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0608_ ) );
MUX2_X1 \myreg/_4870_ ( .A(\myreg/_0331_ ), .B(\myreg/_2177_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0609_ ) );
MUX2_X1 \myreg/_4871_ ( .A(\myreg/_0342_ ), .B(\myreg/_2179_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0610_ ) );
MUX2_X1 \myreg/_4872_ ( .A(\myreg/_0345_ ), .B(\myreg/_2181_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0611_ ) );
MUX2_X1 \myreg/_4873_ ( .A(\myreg/_0346_ ), .B(\myreg/_2183_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0612_ ) );
MUX2_X1 \myreg/_4874_ ( .A(\myreg/_0347_ ), .B(\myreg/_2185_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0613_ ) );
MUX2_X1 \myreg/_4875_ ( .A(\myreg/_0348_ ), .B(\myreg/_2187_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0614_ ) );
MUX2_X1 \myreg/_4876_ ( .A(\myreg/_0349_ ), .B(\myreg/_2189_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0615_ ) );
MUX2_X1 \myreg/_4877_ ( .A(\myreg/_0350_ ), .B(\myreg/_2191_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0616_ ) );
MUX2_X1 \myreg/_4878_ ( .A(\myreg/_0351_ ), .B(\myreg/_2193_ ), .S(\myreg/_2258_ ), .Z(\myreg/_0617_ ) );
BUF_X8 \myreg/_4879_ ( .A(\myreg/_2257_ ), .Z(\myreg/_2259_ ) );
MUX2_X1 \myreg/_4880_ ( .A(\myreg/_0321_ ), .B(\myreg/_2196_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0618_ ) );
MUX2_X1 \myreg/_4881_ ( .A(\myreg/_0322_ ), .B(\myreg/_2199_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0619_ ) );
MUX2_X1 \myreg/_4882_ ( .A(\myreg/_0323_ ), .B(\myreg/_2201_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0620_ ) );
MUX2_X1 \myreg/_4883_ ( .A(\myreg/_0324_ ), .B(\myreg/_2203_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0621_ ) );
MUX2_X1 \myreg/_4884_ ( .A(\myreg/_0325_ ), .B(\myreg/_2205_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0622_ ) );
MUX2_X1 \myreg/_4885_ ( .A(\myreg/_0326_ ), .B(\myreg/_2207_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0623_ ) );
MUX2_X1 \myreg/_4886_ ( .A(\myreg/_0327_ ), .B(\myreg/_2209_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0624_ ) );
MUX2_X1 \myreg/_4887_ ( .A(\myreg/_0328_ ), .B(\myreg/_2211_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0625_ ) );
MUX2_X1 \myreg/_4888_ ( .A(\myreg/_0329_ ), .B(\myreg/_2213_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0626_ ) );
MUX2_X1 \myreg/_4889_ ( .A(\myreg/_0330_ ), .B(\myreg/_2215_ ), .S(\myreg/_2259_ ), .Z(\myreg/_0627_ ) );
BUF_X8 \myreg/_4890_ ( .A(\myreg/_2257_ ), .Z(\myreg/_2260_ ) );
MUX2_X1 \myreg/_4891_ ( .A(\myreg/_0332_ ), .B(\myreg/_2218_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0628_ ) );
MUX2_X1 \myreg/_4892_ ( .A(\myreg/_0333_ ), .B(\myreg/_2221_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0629_ ) );
MUX2_X1 \myreg/_4893_ ( .A(\myreg/_0334_ ), .B(\myreg/_2223_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0630_ ) );
MUX2_X1 \myreg/_4894_ ( .A(\myreg/_0335_ ), .B(\myreg/_2225_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0631_ ) );
MUX2_X1 \myreg/_4895_ ( .A(\myreg/_0336_ ), .B(\myreg/_2227_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0632_ ) );
MUX2_X1 \myreg/_4896_ ( .A(\myreg/_0337_ ), .B(\myreg/_2229_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0633_ ) );
MUX2_X1 \myreg/_4897_ ( .A(\myreg/_0338_ ), .B(\myreg/_2231_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0634_ ) );
MUX2_X1 \myreg/_4898_ ( .A(\myreg/_0339_ ), .B(\myreg/_2233_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0635_ ) );
MUX2_X1 \myreg/_4899_ ( .A(\myreg/_0340_ ), .B(\myreg/_2235_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0636_ ) );
MUX2_X1 \myreg/_4900_ ( .A(\myreg/_0341_ ), .B(\myreg/_2237_ ), .S(\myreg/_2260_ ), .Z(\myreg/_0637_ ) );
MUX2_X1 \myreg/_4901_ ( .A(\myreg/_0343_ ), .B(\myreg/_2239_ ), .S(\myreg/_2257_ ), .Z(\myreg/_0638_ ) );
MUX2_X1 \myreg/_4902_ ( .A(\myreg/_0344_ ), .B(\myreg/_2241_ ), .S(\myreg/_2257_ ), .Z(\myreg/_0639_ ) );
NOR2_X4 \myreg/_4903_ ( .A1(\myreg/_2170_ ), .A2(\myreg/_2246_ ), .ZN(\myreg/_2261_ ) );
BUF_X8 \myreg/_4904_ ( .A(\myreg/_2261_ ), .Z(\myreg/_2262_ ) );
MUX2_X1 \myreg/_4905_ ( .A(\myreg/_0288_ ), .B(\myreg/_2168_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0640_ ) );
MUX2_X1 \myreg/_4906_ ( .A(\myreg/_0299_ ), .B(\myreg/_2177_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0641_ ) );
MUX2_X1 \myreg/_4907_ ( .A(\myreg/_0310_ ), .B(\myreg/_2179_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0642_ ) );
MUX2_X1 \myreg/_4908_ ( .A(\myreg/_0313_ ), .B(\myreg/_2181_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0643_ ) );
MUX2_X1 \myreg/_4909_ ( .A(\myreg/_0314_ ), .B(\myreg/_2183_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0644_ ) );
MUX2_X1 \myreg/_4910_ ( .A(\myreg/_0315_ ), .B(\myreg/_2185_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0645_ ) );
MUX2_X1 \myreg/_4911_ ( .A(\myreg/_0316_ ), .B(\myreg/_2187_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0646_ ) );
MUX2_X1 \myreg/_4912_ ( .A(\myreg/_0317_ ), .B(\myreg/_2189_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0647_ ) );
MUX2_X1 \myreg/_4913_ ( .A(\myreg/_0318_ ), .B(\myreg/_2191_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0648_ ) );
MUX2_X1 \myreg/_4914_ ( .A(\myreg/_0319_ ), .B(\myreg/_2193_ ), .S(\myreg/_2262_ ), .Z(\myreg/_0649_ ) );
BUF_X8 \myreg/_4915_ ( .A(\myreg/_2261_ ), .Z(\myreg/_2263_ ) );
MUX2_X1 \myreg/_4916_ ( .A(\myreg/_0289_ ), .B(\myreg/_2196_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0650_ ) );
MUX2_X1 \myreg/_4917_ ( .A(\myreg/_0290_ ), .B(\myreg/_2199_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0651_ ) );
MUX2_X1 \myreg/_4918_ ( .A(\myreg/_0291_ ), .B(\myreg/_2201_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0652_ ) );
MUX2_X1 \myreg/_4919_ ( .A(\myreg/_0292_ ), .B(\myreg/_2203_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0653_ ) );
MUX2_X1 \myreg/_4920_ ( .A(\myreg/_0293_ ), .B(\myreg/_2205_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0654_ ) );
MUX2_X1 \myreg/_4921_ ( .A(\myreg/_0294_ ), .B(\myreg/_2207_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0655_ ) );
MUX2_X1 \myreg/_4922_ ( .A(\myreg/_0295_ ), .B(\myreg/_2209_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0656_ ) );
MUX2_X1 \myreg/_4923_ ( .A(\myreg/_0296_ ), .B(\myreg/_2211_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0657_ ) );
MUX2_X1 \myreg/_4924_ ( .A(\myreg/_0297_ ), .B(\myreg/_2213_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0658_ ) );
MUX2_X1 \myreg/_4925_ ( .A(\myreg/_0298_ ), .B(\myreg/_2215_ ), .S(\myreg/_2263_ ), .Z(\myreg/_0659_ ) );
BUF_X8 \myreg/_4926_ ( .A(\myreg/_2261_ ), .Z(\myreg/_2264_ ) );
MUX2_X1 \myreg/_4927_ ( .A(\myreg/_0300_ ), .B(\myreg/_2218_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0660_ ) );
MUX2_X1 \myreg/_4928_ ( .A(\myreg/_0301_ ), .B(\myreg/_2221_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0661_ ) );
MUX2_X1 \myreg/_4929_ ( .A(\myreg/_0302_ ), .B(\myreg/_2223_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0662_ ) );
MUX2_X1 \myreg/_4930_ ( .A(\myreg/_0303_ ), .B(\myreg/_2225_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0663_ ) );
MUX2_X1 \myreg/_4931_ ( .A(\myreg/_0304_ ), .B(\myreg/_2227_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0664_ ) );
MUX2_X1 \myreg/_4932_ ( .A(\myreg/_0305_ ), .B(\myreg/_2229_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0665_ ) );
MUX2_X1 \myreg/_4933_ ( .A(\myreg/_0306_ ), .B(\myreg/_2231_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0666_ ) );
MUX2_X1 \myreg/_4934_ ( .A(\myreg/_0307_ ), .B(\myreg/_2233_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0667_ ) );
MUX2_X1 \myreg/_4935_ ( .A(\myreg/_0308_ ), .B(\myreg/_2235_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0668_ ) );
MUX2_X1 \myreg/_4936_ ( .A(\myreg/_0309_ ), .B(\myreg/_2237_ ), .S(\myreg/_2264_ ), .Z(\myreg/_0669_ ) );
MUX2_X1 \myreg/_4937_ ( .A(\myreg/_0311_ ), .B(\myreg/_2239_ ), .S(\myreg/_2261_ ), .Z(\myreg/_0670_ ) );
MUX2_X1 \myreg/_4938_ ( .A(\myreg/_0312_ ), .B(\myreg/_2241_ ), .S(\myreg/_2261_ ), .Z(\myreg/_0671_ ) );
AND2_X4 \myreg/_4939_ ( .A1(\myreg/_2165_ ), .A2(\myreg/_2416_ ), .ZN(\myreg/_2265_ ) );
NAND2_X4 \myreg/_4940_ ( .A1(\myreg/_2265_ ), .A2(\myreg/_2162_ ), .ZN(\myreg/_2266_ ) );
NOR2_X4 \myreg/_4941_ ( .A1(\myreg/_2266_ ), .A2(\myreg/_2256_ ), .ZN(\myreg/_2267_ ) );
BUF_X8 \myreg/_4942_ ( .A(\myreg/_2267_ ), .Z(\myreg/_2268_ ) );
MUX2_X1 \myreg/_4943_ ( .A(\myreg/_0448_ ), .B(\myreg/_2168_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0672_ ) );
MUX2_X1 \myreg/_4944_ ( .A(\myreg/_0459_ ), .B(\myreg/_2177_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0673_ ) );
MUX2_X1 \myreg/_4945_ ( .A(\myreg/_0470_ ), .B(\myreg/_2179_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0674_ ) );
MUX2_X1 \myreg/_4946_ ( .A(\myreg/_0473_ ), .B(\myreg/_2181_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0675_ ) );
MUX2_X1 \myreg/_4947_ ( .A(\myreg/_0474_ ), .B(\myreg/_2183_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0676_ ) );
MUX2_X1 \myreg/_4948_ ( .A(\myreg/_0475_ ), .B(\myreg/_2185_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0677_ ) );
MUX2_X1 \myreg/_4949_ ( .A(\myreg/_0476_ ), .B(\myreg/_2187_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0678_ ) );
MUX2_X1 \myreg/_4950_ ( .A(\myreg/_0477_ ), .B(\myreg/_2189_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0679_ ) );
MUX2_X1 \myreg/_4951_ ( .A(\myreg/_0478_ ), .B(\myreg/_2191_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0680_ ) );
MUX2_X1 \myreg/_4952_ ( .A(\myreg/_0479_ ), .B(\myreg/_2193_ ), .S(\myreg/_2268_ ), .Z(\myreg/_0681_ ) );
BUF_X8 \myreg/_4953_ ( .A(\myreg/_2267_ ), .Z(\myreg/_2269_ ) );
MUX2_X1 \myreg/_4954_ ( .A(\myreg/_0449_ ), .B(\myreg/_2196_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0682_ ) );
MUX2_X1 \myreg/_4955_ ( .A(\myreg/_0450_ ), .B(\myreg/_2199_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0683_ ) );
MUX2_X1 \myreg/_4956_ ( .A(\myreg/_0451_ ), .B(\myreg/_2201_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0684_ ) );
MUX2_X1 \myreg/_4957_ ( .A(\myreg/_0452_ ), .B(\myreg/_2203_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0685_ ) );
MUX2_X1 \myreg/_4958_ ( .A(\myreg/_0453_ ), .B(\myreg/_2205_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0686_ ) );
MUX2_X1 \myreg/_4959_ ( .A(\myreg/_0454_ ), .B(\myreg/_2207_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0687_ ) );
MUX2_X1 \myreg/_4960_ ( .A(\myreg/_0455_ ), .B(\myreg/_2209_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0688_ ) );
MUX2_X1 \myreg/_4961_ ( .A(\myreg/_0456_ ), .B(\myreg/_2211_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0689_ ) );
MUX2_X1 \myreg/_4962_ ( .A(\myreg/_0457_ ), .B(\myreg/_2213_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0690_ ) );
MUX2_X1 \myreg/_4963_ ( .A(\myreg/_0458_ ), .B(\myreg/_2215_ ), .S(\myreg/_2269_ ), .Z(\myreg/_0691_ ) );
BUF_X8 \myreg/_4964_ ( .A(\myreg/_2267_ ), .Z(\myreg/_2270_ ) );
MUX2_X1 \myreg/_4965_ ( .A(\myreg/_0460_ ), .B(\myreg/_2218_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0692_ ) );
MUX2_X1 \myreg/_4966_ ( .A(\myreg/_0461_ ), .B(\myreg/_2221_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0693_ ) );
MUX2_X1 \myreg/_4967_ ( .A(\myreg/_0462_ ), .B(\myreg/_2223_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0694_ ) );
MUX2_X1 \myreg/_4968_ ( .A(\myreg/_0463_ ), .B(\myreg/_2225_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0695_ ) );
MUX2_X1 \myreg/_4969_ ( .A(\myreg/_0464_ ), .B(\myreg/_2227_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0696_ ) );
MUX2_X1 \myreg/_4970_ ( .A(\myreg/_0465_ ), .B(\myreg/_2229_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0697_ ) );
MUX2_X1 \myreg/_4971_ ( .A(\myreg/_0466_ ), .B(\myreg/_2231_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0698_ ) );
MUX2_X1 \myreg/_4972_ ( .A(\myreg/_0467_ ), .B(\myreg/_2233_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0699_ ) );
MUX2_X1 \myreg/_4973_ ( .A(\myreg/_0468_ ), .B(\myreg/_2235_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0700_ ) );
MUX2_X1 \myreg/_4974_ ( .A(\myreg/_0469_ ), .B(\myreg/_2237_ ), .S(\myreg/_2270_ ), .Z(\myreg/_0701_ ) );
MUX2_X1 \myreg/_4975_ ( .A(\myreg/_0471_ ), .B(\myreg/_2239_ ), .S(\myreg/_2267_ ), .Z(\myreg/_0702_ ) );
MUX2_X1 \myreg/_4976_ ( .A(\myreg/_0472_ ), .B(\myreg/_2241_ ), .S(\myreg/_2267_ ), .Z(\myreg/_0703_ ) );
INV_X1 \myreg/_4977_ ( .A(\myreg/_0000_ ), .ZN(\myreg/_2271_ ) );
NOR2_X1 \myreg/_4978_ ( .A1(\myreg/_2271_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0704_ ) );
INV_X1 \myreg/_4979_ ( .A(\myreg/_0011_ ), .ZN(\myreg/_2272_ ) );
NOR2_X1 \myreg/_4980_ ( .A1(\myreg/_2272_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0705_ ) );
INV_X1 \myreg/_4981_ ( .A(\myreg/_0022_ ), .ZN(\myreg/_2273_ ) );
NOR2_X1 \myreg/_4982_ ( .A1(\myreg/_2273_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0706_ ) );
INV_X1 \myreg/_4983_ ( .A(\myreg/_0025_ ), .ZN(\myreg/_2274_ ) );
NOR2_X1 \myreg/_4984_ ( .A1(\myreg/_2274_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0707_ ) );
INV_X1 \myreg/_4985_ ( .A(\myreg/_0026_ ), .ZN(\myreg/_2275_ ) );
NOR2_X1 \myreg/_4986_ ( .A1(\myreg/_2275_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0708_ ) );
INV_X1 \myreg/_4987_ ( .A(\myreg/_0027_ ), .ZN(\myreg/_2276_ ) );
NOR2_X1 \myreg/_4988_ ( .A1(\myreg/_2276_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0709_ ) );
INV_X1 \myreg/_4989_ ( .A(\myreg/_0028_ ), .ZN(\myreg/_2277_ ) );
NOR2_X1 \myreg/_4990_ ( .A1(\myreg/_2277_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0710_ ) );
INV_X1 \myreg/_4991_ ( .A(\myreg/_0029_ ), .ZN(\myreg/_2278_ ) );
NOR2_X1 \myreg/_4992_ ( .A1(\myreg/_2278_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0711_ ) );
INV_X1 \myreg/_4993_ ( .A(\myreg/_0030_ ), .ZN(\myreg/_2279_ ) );
NOR2_X1 \myreg/_4994_ ( .A1(\myreg/_2279_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0712_ ) );
INV_X1 \myreg/_4995_ ( .A(\myreg/_0031_ ), .ZN(\myreg/_2280_ ) );
NOR2_X1 \myreg/_4996_ ( .A1(\myreg/_2280_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0713_ ) );
INV_X1 \myreg/_4997_ ( .A(\myreg/_0001_ ), .ZN(\myreg/_2281_ ) );
NOR2_X1 \myreg/_4998_ ( .A1(\myreg/_2281_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0714_ ) );
INV_X1 \myreg/_4999_ ( .A(\myreg/_0002_ ), .ZN(\myreg/_2282_ ) );
NOR2_X1 \myreg/_5000_ ( .A1(\myreg/_2282_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0715_ ) );
INV_X1 \myreg/_5001_ ( .A(\myreg/_0003_ ), .ZN(\myreg/_2283_ ) );
NOR2_X1 \myreg/_5002_ ( .A1(\myreg/_2283_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0716_ ) );
INV_X1 \myreg/_5003_ ( .A(\myreg/_0004_ ), .ZN(\myreg/_2284_ ) );
NOR2_X1 \myreg/_5004_ ( .A1(\myreg/_2284_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0717_ ) );
INV_X1 \myreg/_5005_ ( .A(\myreg/_0005_ ), .ZN(\myreg/_2285_ ) );
NOR2_X1 \myreg/_5006_ ( .A1(\myreg/_2285_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0718_ ) );
INV_X1 \myreg/_5007_ ( .A(\myreg/_0006_ ), .ZN(\myreg/_2286_ ) );
NOR2_X1 \myreg/_5008_ ( .A1(\myreg/_2286_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0719_ ) );
INV_X1 \myreg/_5009_ ( .A(\myreg/_0007_ ), .ZN(\myreg/_2287_ ) );
NOR2_X1 \myreg/_5010_ ( .A1(\myreg/_2287_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0720_ ) );
INV_X1 \myreg/_5011_ ( .A(\myreg/_0008_ ), .ZN(\myreg/_2288_ ) );
NOR2_X1 \myreg/_5012_ ( .A1(\myreg/_2288_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0721_ ) );
INV_X1 \myreg/_5013_ ( .A(\myreg/_0009_ ), .ZN(\myreg/_2289_ ) );
NOR2_X1 \myreg/_5014_ ( .A1(\myreg/_2289_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0722_ ) );
INV_X1 \myreg/_5015_ ( .A(\myreg/_0010_ ), .ZN(\myreg/_2290_ ) );
NOR2_X1 \myreg/_5016_ ( .A1(\myreg/_2290_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0723_ ) );
INV_X1 \myreg/_5017_ ( .A(\myreg/_0012_ ), .ZN(\myreg/_2291_ ) );
NOR2_X1 \myreg/_5018_ ( .A1(\myreg/_2291_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0724_ ) );
INV_X1 \myreg/_5019_ ( .A(\myreg/_0013_ ), .ZN(\myreg/_2292_ ) );
NOR2_X1 \myreg/_5020_ ( .A1(\myreg/_2292_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0725_ ) );
INV_X1 \myreg/_5021_ ( .A(\myreg/_0014_ ), .ZN(\myreg/_2293_ ) );
NOR2_X1 \myreg/_5022_ ( .A1(\myreg/_2293_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0726_ ) );
INV_X1 \myreg/_5023_ ( .A(\myreg/_0015_ ), .ZN(\myreg/_2294_ ) );
NOR2_X1 \myreg/_5024_ ( .A1(\myreg/_2294_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0727_ ) );
INV_X1 \myreg/_5025_ ( .A(\myreg/_0016_ ), .ZN(\myreg/_2295_ ) );
NOR2_X1 \myreg/_5026_ ( .A1(\myreg/_2295_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0728_ ) );
INV_X1 \myreg/_5027_ ( .A(\myreg/_0017_ ), .ZN(\myreg/_2296_ ) );
NOR2_X1 \myreg/_5028_ ( .A1(\myreg/_2296_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0729_ ) );
INV_X1 \myreg/_5029_ ( .A(\myreg/_0018_ ), .ZN(\myreg/_2297_ ) );
NOR2_X1 \myreg/_5030_ ( .A1(\myreg/_2297_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0730_ ) );
INV_X1 \myreg/_5031_ ( .A(\myreg/_0019_ ), .ZN(\myreg/_2298_ ) );
NOR2_X1 \myreg/_5032_ ( .A1(\myreg/_2298_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0731_ ) );
INV_X1 \myreg/_5033_ ( .A(\myreg/_0020_ ), .ZN(\myreg/_2299_ ) );
NOR2_X1 \myreg/_5034_ ( .A1(\myreg/_2299_ ), .A2(fanout_net_61 ), .ZN(\myreg/_0732_ ) );
INV_X1 \myreg/_5035_ ( .A(\myreg/_0021_ ), .ZN(\myreg/_2300_ ) );
NOR2_X1 \myreg/_5036_ ( .A1(\myreg/_2300_ ), .A2(\myreg/_2412_ ), .ZN(\myreg/_0733_ ) );
INV_X1 \myreg/_5037_ ( .A(\myreg/_0023_ ), .ZN(\myreg/_2301_ ) );
NOR2_X1 \myreg/_5038_ ( .A1(\myreg/_2301_ ), .A2(\myreg/_2412_ ), .ZN(\myreg/_0734_ ) );
INV_X1 \myreg/_5039_ ( .A(\myreg/_0024_ ), .ZN(\myreg/_2302_ ) );
NOR2_X1 \myreg/_5040_ ( .A1(\myreg/_2302_ ), .A2(\myreg/_2412_ ), .ZN(\myreg/_0735_ ) );
NOR2_X4 \myreg/_5041_ ( .A1(\myreg/_2244_ ), .A2(\myreg/_2266_ ), .ZN(\myreg/_2303_ ) );
BUF_X4 \myreg/_5042_ ( .A(\myreg/_2303_ ), .Z(\myreg/_2304_ ) );
MUX2_X1 \myreg/_5043_ ( .A(\myreg/_0032_ ), .B(\myreg/_2168_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0736_ ) );
MUX2_X1 \myreg/_5044_ ( .A(\myreg/_0043_ ), .B(\myreg/_2177_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0737_ ) );
MUX2_X1 \myreg/_5045_ ( .A(\myreg/_0054_ ), .B(\myreg/_2179_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0738_ ) );
MUX2_X1 \myreg/_5046_ ( .A(\myreg/_0057_ ), .B(\myreg/_2181_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0739_ ) );
MUX2_X1 \myreg/_5047_ ( .A(\myreg/_0058_ ), .B(\myreg/_2183_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0740_ ) );
MUX2_X1 \myreg/_5048_ ( .A(\myreg/_0059_ ), .B(\myreg/_2185_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0741_ ) );
MUX2_X1 \myreg/_5049_ ( .A(\myreg/_0060_ ), .B(\myreg/_2187_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0742_ ) );
MUX2_X1 \myreg/_5050_ ( .A(\myreg/_0061_ ), .B(\myreg/_2189_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0743_ ) );
MUX2_X1 \myreg/_5051_ ( .A(\myreg/_0062_ ), .B(\myreg/_2191_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0744_ ) );
MUX2_X1 \myreg/_5052_ ( .A(\myreg/_0063_ ), .B(\myreg/_2193_ ), .S(\myreg/_2304_ ), .Z(\myreg/_0745_ ) );
BUF_X4 \myreg/_5053_ ( .A(\myreg/_2303_ ), .Z(\myreg/_2305_ ) );
MUX2_X1 \myreg/_5054_ ( .A(\myreg/_0033_ ), .B(\myreg/_2196_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0746_ ) );
MUX2_X1 \myreg/_5055_ ( .A(\myreg/_0034_ ), .B(\myreg/_2199_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0747_ ) );
MUX2_X1 \myreg/_5056_ ( .A(\myreg/_0035_ ), .B(\myreg/_2201_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0748_ ) );
MUX2_X1 \myreg/_5057_ ( .A(\myreg/_0036_ ), .B(\myreg/_2203_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0749_ ) );
MUX2_X1 \myreg/_5058_ ( .A(\myreg/_0037_ ), .B(\myreg/_2205_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0750_ ) );
MUX2_X1 \myreg/_5059_ ( .A(\myreg/_0038_ ), .B(\myreg/_2207_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0751_ ) );
MUX2_X1 \myreg/_5060_ ( .A(\myreg/_0039_ ), .B(\myreg/_2209_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0752_ ) );
MUX2_X1 \myreg/_5061_ ( .A(\myreg/_0040_ ), .B(\myreg/_2211_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0753_ ) );
MUX2_X1 \myreg/_5062_ ( .A(\myreg/_0041_ ), .B(\myreg/_2213_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0754_ ) );
MUX2_X1 \myreg/_5063_ ( .A(\myreg/_0042_ ), .B(\myreg/_2215_ ), .S(\myreg/_2305_ ), .Z(\myreg/_0755_ ) );
BUF_X4 \myreg/_5064_ ( .A(\myreg/_2303_ ), .Z(\myreg/_2306_ ) );
MUX2_X1 \myreg/_5065_ ( .A(\myreg/_0044_ ), .B(\myreg/_2218_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0756_ ) );
MUX2_X1 \myreg/_5066_ ( .A(\myreg/_0045_ ), .B(\myreg/_2221_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0757_ ) );
MUX2_X1 \myreg/_5067_ ( .A(\myreg/_0046_ ), .B(\myreg/_2223_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0758_ ) );
MUX2_X1 \myreg/_5068_ ( .A(\myreg/_0047_ ), .B(\myreg/_2225_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0759_ ) );
MUX2_X1 \myreg/_5069_ ( .A(\myreg/_0048_ ), .B(\myreg/_2227_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0760_ ) );
MUX2_X1 \myreg/_5070_ ( .A(\myreg/_0049_ ), .B(\myreg/_2229_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0761_ ) );
MUX2_X1 \myreg/_5071_ ( .A(\myreg/_0050_ ), .B(\myreg/_2231_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0762_ ) );
MUX2_X1 \myreg/_5072_ ( .A(\myreg/_0051_ ), .B(\myreg/_2233_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0763_ ) );
MUX2_X1 \myreg/_5073_ ( .A(\myreg/_0052_ ), .B(\myreg/_2235_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0764_ ) );
MUX2_X1 \myreg/_5074_ ( .A(\myreg/_0053_ ), .B(\myreg/_2237_ ), .S(\myreg/_2306_ ), .Z(\myreg/_0765_ ) );
MUX2_X1 \myreg/_5075_ ( .A(\myreg/_0055_ ), .B(\myreg/_2239_ ), .S(\myreg/_2303_ ), .Z(\myreg/_0766_ ) );
MUX2_X1 \myreg/_5076_ ( .A(\myreg/_0056_ ), .B(\myreg/_2241_ ), .S(\myreg/_2303_ ), .Z(\myreg/_0767_ ) );
NOR2_X4 \myreg/_5077_ ( .A1(\myreg/_2170_ ), .A2(\myreg/_2266_ ), .ZN(\myreg/_2307_ ) );
BUF_X4 \myreg/_5078_ ( .A(\myreg/_2307_ ), .Z(\myreg/_2308_ ) );
MUX2_X1 \myreg/_5079_ ( .A(\myreg/_0064_ ), .B(\myreg/_2168_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0768_ ) );
MUX2_X1 \myreg/_5080_ ( .A(\myreg/_0075_ ), .B(\myreg/_2177_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0769_ ) );
MUX2_X1 \myreg/_5081_ ( .A(\myreg/_0086_ ), .B(\myreg/_2179_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0770_ ) );
MUX2_X1 \myreg/_5082_ ( .A(\myreg/_0089_ ), .B(\myreg/_2181_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0771_ ) );
MUX2_X1 \myreg/_5083_ ( .A(\myreg/_0090_ ), .B(\myreg/_2183_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0772_ ) );
MUX2_X1 \myreg/_5084_ ( .A(\myreg/_0091_ ), .B(\myreg/_2185_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0773_ ) );
MUX2_X1 \myreg/_5085_ ( .A(\myreg/_0092_ ), .B(\myreg/_2187_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0774_ ) );
MUX2_X1 \myreg/_5086_ ( .A(\myreg/_0093_ ), .B(\myreg/_2189_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0775_ ) );
MUX2_X1 \myreg/_5087_ ( .A(\myreg/_0094_ ), .B(\myreg/_2191_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0776_ ) );
MUX2_X1 \myreg/_5088_ ( .A(\myreg/_0095_ ), .B(\myreg/_2193_ ), .S(\myreg/_2308_ ), .Z(\myreg/_0777_ ) );
BUF_X4 \myreg/_5089_ ( .A(\myreg/_2307_ ), .Z(\myreg/_2309_ ) );
MUX2_X1 \myreg/_5090_ ( .A(\myreg/_0065_ ), .B(\myreg/_2196_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0778_ ) );
MUX2_X1 \myreg/_5091_ ( .A(\myreg/_0066_ ), .B(\myreg/_2199_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0779_ ) );
MUX2_X1 \myreg/_5092_ ( .A(\myreg/_0067_ ), .B(\myreg/_2201_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0780_ ) );
MUX2_X1 \myreg/_5093_ ( .A(\myreg/_0068_ ), .B(\myreg/_2203_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0781_ ) );
MUX2_X1 \myreg/_5094_ ( .A(\myreg/_0069_ ), .B(\myreg/_2205_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0782_ ) );
MUX2_X1 \myreg/_5095_ ( .A(\myreg/_0070_ ), .B(\myreg/_2207_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0783_ ) );
MUX2_X1 \myreg/_5096_ ( .A(\myreg/_0071_ ), .B(\myreg/_2209_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0784_ ) );
MUX2_X1 \myreg/_5097_ ( .A(\myreg/_0072_ ), .B(\myreg/_2211_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0785_ ) );
MUX2_X1 \myreg/_5098_ ( .A(\myreg/_0073_ ), .B(\myreg/_2213_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0786_ ) );
MUX2_X1 \myreg/_5099_ ( .A(\myreg/_0074_ ), .B(\myreg/_2215_ ), .S(\myreg/_2309_ ), .Z(\myreg/_0787_ ) );
BUF_X4 \myreg/_5100_ ( .A(\myreg/_2307_ ), .Z(\myreg/_2310_ ) );
MUX2_X1 \myreg/_5101_ ( .A(\myreg/_0076_ ), .B(\myreg/_2218_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0788_ ) );
MUX2_X1 \myreg/_5102_ ( .A(\myreg/_0077_ ), .B(\myreg/_2221_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0789_ ) );
MUX2_X1 \myreg/_5103_ ( .A(\myreg/_0078_ ), .B(\myreg/_2223_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0790_ ) );
MUX2_X1 \myreg/_5104_ ( .A(\myreg/_0079_ ), .B(\myreg/_2225_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0791_ ) );
MUX2_X1 \myreg/_5105_ ( .A(\myreg/_0080_ ), .B(\myreg/_2227_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0792_ ) );
MUX2_X1 \myreg/_5106_ ( .A(\myreg/_0081_ ), .B(\myreg/_2229_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0793_ ) );
MUX2_X1 \myreg/_5107_ ( .A(\myreg/_0082_ ), .B(\myreg/_2231_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0794_ ) );
MUX2_X1 \myreg/_5108_ ( .A(\myreg/_0083_ ), .B(\myreg/_2233_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0795_ ) );
MUX2_X1 \myreg/_5109_ ( .A(\myreg/_0084_ ), .B(\myreg/_2235_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0796_ ) );
MUX2_X1 \myreg/_5110_ ( .A(\myreg/_0085_ ), .B(\myreg/_2237_ ), .S(\myreg/_2310_ ), .Z(\myreg/_0797_ ) );
MUX2_X1 \myreg/_5111_ ( .A(\myreg/_0087_ ), .B(\myreg/_2239_ ), .S(\myreg/_2307_ ), .Z(\myreg/_0798_ ) );
MUX2_X1 \myreg/_5112_ ( .A(\myreg/_0088_ ), .B(\myreg/_2241_ ), .S(\myreg/_2307_ ), .Z(\myreg/_0799_ ) );
NAND2_X4 \myreg/_5113_ ( .A1(\myreg/_2171_ ), .A2(\myreg/_2416_ ), .ZN(\myreg/_2311_ ) );
NOR2_X4 \myreg/_5114_ ( .A1(\myreg/_2311_ ), .A2(\myreg/_2256_ ), .ZN(\myreg/_2312_ ) );
BUF_X8 \myreg/_5115_ ( .A(\myreg/_2312_ ), .Z(\myreg/_2313_ ) );
MUX2_X1 \myreg/_5116_ ( .A(\myreg/_0096_ ), .B(\myreg/_2168_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0800_ ) );
MUX2_X1 \myreg/_5117_ ( .A(\myreg/_0107_ ), .B(\myreg/_2177_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0801_ ) );
MUX2_X1 \myreg/_5118_ ( .A(\myreg/_0118_ ), .B(\myreg/_2179_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0802_ ) );
MUX2_X1 \myreg/_5119_ ( .A(\myreg/_0121_ ), .B(\myreg/_2181_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0803_ ) );
MUX2_X1 \myreg/_5120_ ( .A(\myreg/_0122_ ), .B(\myreg/_2183_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0804_ ) );
MUX2_X1 \myreg/_5121_ ( .A(\myreg/_0123_ ), .B(\myreg/_2185_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0805_ ) );
MUX2_X1 \myreg/_5122_ ( .A(\myreg/_0124_ ), .B(\myreg/_2187_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0806_ ) );
MUX2_X1 \myreg/_5123_ ( .A(\myreg/_0125_ ), .B(\myreg/_2189_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0807_ ) );
MUX2_X1 \myreg/_5124_ ( .A(\myreg/_0126_ ), .B(\myreg/_2191_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0808_ ) );
MUX2_X1 \myreg/_5125_ ( .A(\myreg/_0127_ ), .B(\myreg/_2193_ ), .S(\myreg/_2313_ ), .Z(\myreg/_0809_ ) );
BUF_X8 \myreg/_5126_ ( .A(\myreg/_2312_ ), .Z(\myreg/_2314_ ) );
MUX2_X1 \myreg/_5127_ ( .A(\myreg/_0097_ ), .B(\myreg/_2196_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0810_ ) );
MUX2_X1 \myreg/_5128_ ( .A(\myreg/_0098_ ), .B(\myreg/_2199_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0811_ ) );
MUX2_X1 \myreg/_5129_ ( .A(\myreg/_0099_ ), .B(\myreg/_2201_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0812_ ) );
MUX2_X1 \myreg/_5130_ ( .A(\myreg/_0100_ ), .B(\myreg/_2203_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0813_ ) );
MUX2_X1 \myreg/_5131_ ( .A(\myreg/_0101_ ), .B(\myreg/_2205_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0814_ ) );
MUX2_X1 \myreg/_5132_ ( .A(\myreg/_0102_ ), .B(\myreg/_2207_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0815_ ) );
MUX2_X1 \myreg/_5133_ ( .A(\myreg/_0103_ ), .B(\myreg/_2209_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0816_ ) );
MUX2_X1 \myreg/_5134_ ( .A(\myreg/_0104_ ), .B(\myreg/_2211_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0817_ ) );
MUX2_X1 \myreg/_5135_ ( .A(\myreg/_0105_ ), .B(\myreg/_2213_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0818_ ) );
MUX2_X1 \myreg/_5136_ ( .A(\myreg/_0106_ ), .B(\myreg/_2215_ ), .S(\myreg/_2314_ ), .Z(\myreg/_0819_ ) );
BUF_X8 \myreg/_5137_ ( .A(\myreg/_2312_ ), .Z(\myreg/_2315_ ) );
MUX2_X1 \myreg/_5138_ ( .A(\myreg/_0108_ ), .B(\myreg/_2218_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0820_ ) );
MUX2_X1 \myreg/_5139_ ( .A(\myreg/_0109_ ), .B(\myreg/_2221_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0821_ ) );
MUX2_X1 \myreg/_5140_ ( .A(\myreg/_0110_ ), .B(\myreg/_2223_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0822_ ) );
MUX2_X1 \myreg/_5141_ ( .A(\myreg/_0111_ ), .B(\myreg/_2225_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0823_ ) );
MUX2_X1 \myreg/_5142_ ( .A(\myreg/_0112_ ), .B(\myreg/_2227_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0824_ ) );
MUX2_X1 \myreg/_5143_ ( .A(\myreg/_0113_ ), .B(\myreg/_2229_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0825_ ) );
MUX2_X1 \myreg/_5144_ ( .A(\myreg/_0114_ ), .B(\myreg/_2231_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0826_ ) );
MUX2_X1 \myreg/_5145_ ( .A(\myreg/_0115_ ), .B(\myreg/_2233_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0827_ ) );
MUX2_X1 \myreg/_5146_ ( .A(\myreg/_0116_ ), .B(\myreg/_2235_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0828_ ) );
MUX2_X1 \myreg/_5147_ ( .A(\myreg/_0117_ ), .B(\myreg/_2237_ ), .S(\myreg/_2315_ ), .Z(\myreg/_0829_ ) );
MUX2_X1 \myreg/_5148_ ( .A(\myreg/_0119_ ), .B(\myreg/_2239_ ), .S(\myreg/_2312_ ), .Z(\myreg/_0830_ ) );
MUX2_X1 \myreg/_5149_ ( .A(\myreg/_0120_ ), .B(\myreg/_2241_ ), .S(\myreg/_2312_ ), .Z(\myreg/_0831_ ) );
NOR2_X4 \myreg/_5150_ ( .A1(\myreg/_2251_ ), .A2(\myreg/_2311_ ), .ZN(\myreg/_2316_ ) );
BUF_X4 \myreg/_5151_ ( .A(\myreg/_2316_ ), .Z(\myreg/_2317_ ) );
MUX2_X1 \myreg/_5152_ ( .A(\myreg/_0128_ ), .B(\myreg/_2168_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0832_ ) );
MUX2_X1 \myreg/_5153_ ( .A(\myreg/_0139_ ), .B(\myreg/_2177_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0833_ ) );
MUX2_X1 \myreg/_5154_ ( .A(\myreg/_0150_ ), .B(\myreg/_2179_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0834_ ) );
MUX2_X1 \myreg/_5155_ ( .A(\myreg/_0153_ ), .B(\myreg/_2181_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0835_ ) );
MUX2_X1 \myreg/_5156_ ( .A(\myreg/_0154_ ), .B(\myreg/_2183_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0836_ ) );
MUX2_X1 \myreg/_5157_ ( .A(\myreg/_0155_ ), .B(\myreg/_2185_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0837_ ) );
MUX2_X1 \myreg/_5158_ ( .A(\myreg/_0156_ ), .B(\myreg/_2187_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0838_ ) );
MUX2_X1 \myreg/_5159_ ( .A(\myreg/_0157_ ), .B(\myreg/_2189_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0839_ ) );
MUX2_X1 \myreg/_5160_ ( .A(\myreg/_0158_ ), .B(\myreg/_2191_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0840_ ) );
MUX2_X1 \myreg/_5161_ ( .A(\myreg/_0159_ ), .B(\myreg/_2193_ ), .S(\myreg/_2317_ ), .Z(\myreg/_0841_ ) );
BUF_X4 \myreg/_5162_ ( .A(\myreg/_2316_ ), .Z(\myreg/_2318_ ) );
MUX2_X1 \myreg/_5163_ ( .A(\myreg/_0129_ ), .B(\myreg/_2196_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0842_ ) );
MUX2_X1 \myreg/_5164_ ( .A(\myreg/_0130_ ), .B(\myreg/_2199_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0843_ ) );
MUX2_X1 \myreg/_5165_ ( .A(\myreg/_0131_ ), .B(\myreg/_2201_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0844_ ) );
MUX2_X1 \myreg/_5166_ ( .A(\myreg/_0132_ ), .B(\myreg/_2203_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0845_ ) );
MUX2_X1 \myreg/_5167_ ( .A(\myreg/_0133_ ), .B(\myreg/_2205_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0846_ ) );
MUX2_X1 \myreg/_5168_ ( .A(\myreg/_0134_ ), .B(\myreg/_2207_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0847_ ) );
MUX2_X1 \myreg/_5169_ ( .A(\myreg/_0135_ ), .B(\myreg/_2209_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0848_ ) );
MUX2_X1 \myreg/_5170_ ( .A(\myreg/_0136_ ), .B(\myreg/_2211_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0849_ ) );
MUX2_X1 \myreg/_5171_ ( .A(\myreg/_0137_ ), .B(\myreg/_2213_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0850_ ) );
MUX2_X1 \myreg/_5172_ ( .A(\myreg/_0138_ ), .B(\myreg/_2215_ ), .S(\myreg/_2318_ ), .Z(\myreg/_0851_ ) );
BUF_X4 \myreg/_5173_ ( .A(\myreg/_2316_ ), .Z(\myreg/_2319_ ) );
MUX2_X1 \myreg/_5174_ ( .A(\myreg/_0140_ ), .B(\myreg/_2218_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0852_ ) );
MUX2_X1 \myreg/_5175_ ( .A(\myreg/_0141_ ), .B(\myreg/_2221_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0853_ ) );
MUX2_X1 \myreg/_5176_ ( .A(\myreg/_0142_ ), .B(\myreg/_2223_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0854_ ) );
MUX2_X1 \myreg/_5177_ ( .A(\myreg/_0143_ ), .B(\myreg/_2225_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0855_ ) );
MUX2_X1 \myreg/_5178_ ( .A(\myreg/_0144_ ), .B(\myreg/_2227_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0856_ ) );
MUX2_X1 \myreg/_5179_ ( .A(\myreg/_0145_ ), .B(\myreg/_2229_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0857_ ) );
MUX2_X1 \myreg/_5180_ ( .A(\myreg/_0146_ ), .B(\myreg/_2231_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0858_ ) );
MUX2_X1 \myreg/_5181_ ( .A(\myreg/_0147_ ), .B(\myreg/_2233_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0859_ ) );
MUX2_X1 \myreg/_5182_ ( .A(\myreg/_0148_ ), .B(\myreg/_2235_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0860_ ) );
MUX2_X1 \myreg/_5183_ ( .A(\myreg/_0149_ ), .B(\myreg/_2237_ ), .S(\myreg/_2319_ ), .Z(\myreg/_0861_ ) );
MUX2_X1 \myreg/_5184_ ( .A(\myreg/_0151_ ), .B(\myreg/_2239_ ), .S(\myreg/_2316_ ), .Z(\myreg/_0862_ ) );
MUX2_X1 \myreg/_5185_ ( .A(\myreg/_0152_ ), .B(\myreg/_2241_ ), .S(\myreg/_2316_ ), .Z(\myreg/_0863_ ) );
NOR2_X4 \myreg/_5186_ ( .A1(\myreg/_2244_ ), .A2(\myreg/_2311_ ), .ZN(\myreg/_2320_ ) );
BUF_X4 \myreg/_5187_ ( .A(\myreg/_2320_ ), .Z(\myreg/_2321_ ) );
MUX2_X1 \myreg/_5188_ ( .A(\myreg/_0160_ ), .B(\myreg/_2167_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0864_ ) );
MUX2_X1 \myreg/_5189_ ( .A(\myreg/_0171_ ), .B(\myreg/_2176_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0865_ ) );
MUX2_X1 \myreg/_5190_ ( .A(\myreg/_0182_ ), .B(\myreg/_2178_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0866_ ) );
MUX2_X1 \myreg/_5191_ ( .A(\myreg/_0185_ ), .B(\myreg/_2180_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0867_ ) );
MUX2_X1 \myreg/_5192_ ( .A(\myreg/_0186_ ), .B(\myreg/_2182_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0868_ ) );
MUX2_X1 \myreg/_5193_ ( .A(\myreg/_0187_ ), .B(\myreg/_2184_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0869_ ) );
MUX2_X1 \myreg/_5194_ ( .A(\myreg/_0188_ ), .B(\myreg/_2186_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0870_ ) );
MUX2_X1 \myreg/_5195_ ( .A(\myreg/_0189_ ), .B(\myreg/_2188_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0871_ ) );
MUX2_X1 \myreg/_5196_ ( .A(\myreg/_0190_ ), .B(\myreg/_2190_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0872_ ) );
MUX2_X1 \myreg/_5197_ ( .A(\myreg/_0191_ ), .B(\myreg/_2192_ ), .S(\myreg/_2321_ ), .Z(\myreg/_0873_ ) );
BUF_X4 \myreg/_5198_ ( .A(\myreg/_2320_ ), .Z(\myreg/_2322_ ) );
MUX2_X1 \myreg/_5199_ ( .A(\myreg/_0161_ ), .B(\myreg/_2195_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0874_ ) );
MUX2_X1 \myreg/_5200_ ( .A(\myreg/_0162_ ), .B(\myreg/_2198_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0875_ ) );
MUX2_X1 \myreg/_5201_ ( .A(\myreg/_0163_ ), .B(\myreg/_2200_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0876_ ) );
MUX2_X1 \myreg/_5202_ ( .A(\myreg/_0164_ ), .B(\myreg/_2202_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0877_ ) );
MUX2_X1 \myreg/_5203_ ( .A(\myreg/_0165_ ), .B(\myreg/_2204_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0878_ ) );
MUX2_X1 \myreg/_5204_ ( .A(\myreg/_0166_ ), .B(\myreg/_2206_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0879_ ) );
MUX2_X1 \myreg/_5205_ ( .A(\myreg/_0167_ ), .B(\myreg/_2208_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0880_ ) );
MUX2_X1 \myreg/_5206_ ( .A(\myreg/_0168_ ), .B(\myreg/_2210_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0881_ ) );
MUX2_X1 \myreg/_5207_ ( .A(\myreg/_0169_ ), .B(\myreg/_2212_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0882_ ) );
MUX2_X1 \myreg/_5208_ ( .A(\myreg/_0170_ ), .B(\myreg/_2214_ ), .S(\myreg/_2322_ ), .Z(\myreg/_0883_ ) );
BUF_X4 \myreg/_5209_ ( .A(\myreg/_2320_ ), .Z(\myreg/_2323_ ) );
MUX2_X1 \myreg/_5210_ ( .A(\myreg/_0172_ ), .B(\myreg/_2217_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0884_ ) );
MUX2_X1 \myreg/_5211_ ( .A(\myreg/_0173_ ), .B(\myreg/_2220_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0885_ ) );
MUX2_X1 \myreg/_5212_ ( .A(\myreg/_0174_ ), .B(\myreg/_2222_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0886_ ) );
MUX2_X1 \myreg/_5213_ ( .A(\myreg/_0175_ ), .B(\myreg/_2224_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0887_ ) );
MUX2_X1 \myreg/_5214_ ( .A(\myreg/_0176_ ), .B(\myreg/_2226_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0888_ ) );
MUX2_X1 \myreg/_5215_ ( .A(\myreg/_0177_ ), .B(\myreg/_2228_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0889_ ) );
MUX2_X1 \myreg/_5216_ ( .A(\myreg/_0178_ ), .B(\myreg/_2230_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0890_ ) );
MUX2_X1 \myreg/_5217_ ( .A(\myreg/_0179_ ), .B(\myreg/_2232_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0891_ ) );
MUX2_X1 \myreg/_5218_ ( .A(\myreg/_0180_ ), .B(\myreg/_2234_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0892_ ) );
MUX2_X1 \myreg/_5219_ ( .A(\myreg/_0181_ ), .B(\myreg/_2236_ ), .S(\myreg/_2323_ ), .Z(\myreg/_0893_ ) );
MUX2_X1 \myreg/_5220_ ( .A(\myreg/_0183_ ), .B(\myreg/_2238_ ), .S(\myreg/_2320_ ), .Z(\myreg/_0894_ ) );
MUX2_X1 \myreg/_5221_ ( .A(\myreg/_0184_ ), .B(\myreg/_2240_ ), .S(\myreg/_2320_ ), .Z(\myreg/_0895_ ) );
NOR2_X4 \myreg/_5222_ ( .A1(\myreg/_2173_ ), .A2(\myreg/_2244_ ), .ZN(\myreg/_2324_ ) );
BUF_X4 \myreg/_5223_ ( .A(\myreg/_2324_ ), .Z(\myreg/_2325_ ) );
MUX2_X1 \myreg/_5224_ ( .A(\myreg/_0384_ ), .B(\myreg/_2167_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0896_ ) );
MUX2_X1 \myreg/_5225_ ( .A(\myreg/_0395_ ), .B(\myreg/_2176_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0897_ ) );
MUX2_X1 \myreg/_5226_ ( .A(\myreg/_0406_ ), .B(\myreg/_2178_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0898_ ) );
MUX2_X1 \myreg/_5227_ ( .A(\myreg/_0409_ ), .B(\myreg/_2180_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0899_ ) );
MUX2_X1 \myreg/_5228_ ( .A(\myreg/_0410_ ), .B(\myreg/_2182_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0900_ ) );
MUX2_X1 \myreg/_5229_ ( .A(\myreg/_0411_ ), .B(\myreg/_2184_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0901_ ) );
MUX2_X1 \myreg/_5230_ ( .A(\myreg/_0412_ ), .B(\myreg/_2186_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0902_ ) );
MUX2_X1 \myreg/_5231_ ( .A(\myreg/_0413_ ), .B(\myreg/_2188_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0903_ ) );
MUX2_X1 \myreg/_5232_ ( .A(\myreg/_0414_ ), .B(\myreg/_2190_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0904_ ) );
MUX2_X1 \myreg/_5233_ ( .A(\myreg/_0415_ ), .B(\myreg/_2192_ ), .S(\myreg/_2325_ ), .Z(\myreg/_0905_ ) );
BUF_X4 \myreg/_5234_ ( .A(\myreg/_2324_ ), .Z(\myreg/_2326_ ) );
MUX2_X1 \myreg/_5235_ ( .A(\myreg/_0385_ ), .B(\myreg/_2195_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0906_ ) );
MUX2_X1 \myreg/_5236_ ( .A(\myreg/_0386_ ), .B(\myreg/_2198_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0907_ ) );
MUX2_X1 \myreg/_5237_ ( .A(\myreg/_0387_ ), .B(\myreg/_2200_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0908_ ) );
MUX2_X1 \myreg/_5238_ ( .A(\myreg/_0388_ ), .B(\myreg/_2202_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0909_ ) );
MUX2_X1 \myreg/_5239_ ( .A(\myreg/_0389_ ), .B(\myreg/_2204_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0910_ ) );
MUX2_X1 \myreg/_5240_ ( .A(\myreg/_0390_ ), .B(\myreg/_2206_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0911_ ) );
MUX2_X1 \myreg/_5241_ ( .A(\myreg/_0391_ ), .B(\myreg/_2208_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0912_ ) );
MUX2_X1 \myreg/_5242_ ( .A(\myreg/_0392_ ), .B(\myreg/_2210_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0913_ ) );
MUX2_X1 \myreg/_5243_ ( .A(\myreg/_0393_ ), .B(\myreg/_2212_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0914_ ) );
MUX2_X1 \myreg/_5244_ ( .A(\myreg/_0394_ ), .B(\myreg/_2214_ ), .S(\myreg/_2326_ ), .Z(\myreg/_0915_ ) );
BUF_X4 \myreg/_5245_ ( .A(\myreg/_2324_ ), .Z(\myreg/_2327_ ) );
MUX2_X1 \myreg/_5246_ ( .A(\myreg/_0396_ ), .B(\myreg/_2217_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0916_ ) );
MUX2_X1 \myreg/_5247_ ( .A(\myreg/_0397_ ), .B(\myreg/_2220_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0917_ ) );
MUX2_X1 \myreg/_5248_ ( .A(\myreg/_0398_ ), .B(\myreg/_2222_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0918_ ) );
MUX2_X1 \myreg/_5249_ ( .A(\myreg/_0399_ ), .B(\myreg/_2224_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0919_ ) );
MUX2_X1 \myreg/_5250_ ( .A(\myreg/_0400_ ), .B(\myreg/_2226_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0920_ ) );
MUX2_X1 \myreg/_5251_ ( .A(\myreg/_0401_ ), .B(\myreg/_2228_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0921_ ) );
MUX2_X1 \myreg/_5252_ ( .A(\myreg/_0402_ ), .B(\myreg/_2230_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0922_ ) );
MUX2_X1 \myreg/_5253_ ( .A(\myreg/_0403_ ), .B(\myreg/_2232_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0923_ ) );
MUX2_X1 \myreg/_5254_ ( .A(\myreg/_0404_ ), .B(\myreg/_2234_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0924_ ) );
MUX2_X1 \myreg/_5255_ ( .A(\myreg/_0405_ ), .B(\myreg/_2236_ ), .S(\myreg/_2327_ ), .Z(\myreg/_0925_ ) );
MUX2_X1 \myreg/_5256_ ( .A(\myreg/_0407_ ), .B(\myreg/_2238_ ), .S(\myreg/_2324_ ), .Z(\myreg/_0926_ ) );
MUX2_X1 \myreg/_5257_ ( .A(\myreg/_0408_ ), .B(\myreg/_2240_ ), .S(\myreg/_2324_ ), .Z(\myreg/_0927_ ) );
NOR2_X4 \myreg/_5258_ ( .A1(\myreg/_2170_ ), .A2(\myreg/_2311_ ), .ZN(\myreg/_2328_ ) );
BUF_X4 \myreg/_5259_ ( .A(\myreg/_2328_ ), .Z(\myreg/_2329_ ) );
MUX2_X1 \myreg/_5260_ ( .A(\myreg/_0192_ ), .B(\myreg/_2167_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0928_ ) );
MUX2_X1 \myreg/_5261_ ( .A(\myreg/_0203_ ), .B(\myreg/_2176_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0929_ ) );
MUX2_X1 \myreg/_5262_ ( .A(\myreg/_0214_ ), .B(\myreg/_2178_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0930_ ) );
MUX2_X1 \myreg/_5263_ ( .A(\myreg/_0217_ ), .B(\myreg/_2180_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0931_ ) );
MUX2_X1 \myreg/_5264_ ( .A(\myreg/_0218_ ), .B(\myreg/_2182_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0932_ ) );
MUX2_X1 \myreg/_5265_ ( .A(\myreg/_0219_ ), .B(\myreg/_2184_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0933_ ) );
MUX2_X1 \myreg/_5266_ ( .A(\myreg/_0220_ ), .B(\myreg/_2186_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0934_ ) );
MUX2_X1 \myreg/_5267_ ( .A(\myreg/_0221_ ), .B(\myreg/_2188_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0935_ ) );
MUX2_X1 \myreg/_5268_ ( .A(\myreg/_0222_ ), .B(\myreg/_2190_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0936_ ) );
MUX2_X1 \myreg/_5269_ ( .A(\myreg/_0223_ ), .B(\myreg/_2192_ ), .S(\myreg/_2329_ ), .Z(\myreg/_0937_ ) );
BUF_X4 \myreg/_5270_ ( .A(\myreg/_2328_ ), .Z(\myreg/_2330_ ) );
MUX2_X1 \myreg/_5271_ ( .A(\myreg/_0193_ ), .B(\myreg/_2195_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0938_ ) );
MUX2_X1 \myreg/_5272_ ( .A(\myreg/_0194_ ), .B(\myreg/_2198_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0939_ ) );
MUX2_X1 \myreg/_5273_ ( .A(\myreg/_0195_ ), .B(\myreg/_2200_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0940_ ) );
MUX2_X1 \myreg/_5274_ ( .A(\myreg/_0196_ ), .B(\myreg/_2202_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0941_ ) );
MUX2_X1 \myreg/_5275_ ( .A(\myreg/_0197_ ), .B(\myreg/_2204_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0942_ ) );
MUX2_X1 \myreg/_5276_ ( .A(\myreg/_0198_ ), .B(\myreg/_2206_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0943_ ) );
MUX2_X1 \myreg/_5277_ ( .A(\myreg/_0199_ ), .B(\myreg/_2208_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0944_ ) );
MUX2_X1 \myreg/_5278_ ( .A(\myreg/_0200_ ), .B(\myreg/_2210_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0945_ ) );
MUX2_X1 \myreg/_5279_ ( .A(\myreg/_0201_ ), .B(\myreg/_2212_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0946_ ) );
MUX2_X1 \myreg/_5280_ ( .A(\myreg/_0202_ ), .B(\myreg/_2214_ ), .S(\myreg/_2330_ ), .Z(\myreg/_0947_ ) );
BUF_X4 \myreg/_5281_ ( .A(\myreg/_2328_ ), .Z(\myreg/_2331_ ) );
MUX2_X1 \myreg/_5282_ ( .A(\myreg/_0204_ ), .B(\myreg/_2217_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0948_ ) );
MUX2_X1 \myreg/_5283_ ( .A(\myreg/_0205_ ), .B(\myreg/_2220_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0949_ ) );
MUX2_X1 \myreg/_5284_ ( .A(\myreg/_0206_ ), .B(\myreg/_2222_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0950_ ) );
MUX2_X1 \myreg/_5285_ ( .A(\myreg/_0207_ ), .B(\myreg/_2224_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0951_ ) );
MUX2_X1 \myreg/_5286_ ( .A(\myreg/_0208_ ), .B(\myreg/_2226_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0952_ ) );
MUX2_X1 \myreg/_5287_ ( .A(\myreg/_0209_ ), .B(\myreg/_2228_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0953_ ) );
MUX2_X1 \myreg/_5288_ ( .A(\myreg/_0210_ ), .B(\myreg/_2230_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0954_ ) );
MUX2_X1 \myreg/_5289_ ( .A(\myreg/_0211_ ), .B(\myreg/_2232_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0955_ ) );
MUX2_X1 \myreg/_5290_ ( .A(\myreg/_0212_ ), .B(\myreg/_2234_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0956_ ) );
MUX2_X1 \myreg/_5291_ ( .A(\myreg/_0213_ ), .B(\myreg/_2236_ ), .S(\myreg/_2331_ ), .Z(\myreg/_0957_ ) );
MUX2_X1 \myreg/_5292_ ( .A(\myreg/_0215_ ), .B(\myreg/_2238_ ), .S(\myreg/_2328_ ), .Z(\myreg/_0958_ ) );
MUX2_X1 \myreg/_5293_ ( .A(\myreg/_0216_ ), .B(\myreg/_2240_ ), .S(\myreg/_2328_ ), .Z(\myreg/_0959_ ) );
NOR2_X4 \myreg/_5294_ ( .A1(\myreg/_2251_ ), .A2(\myreg/_2266_ ), .ZN(\myreg/_2332_ ) );
BUF_X4 \myreg/_5295_ ( .A(\myreg/_2332_ ), .Z(\myreg/_2333_ ) );
MUX2_X1 \myreg/_5296_ ( .A(\myreg/_0480_ ), .B(\myreg/_2167_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0960_ ) );
MUX2_X1 \myreg/_5297_ ( .A(\myreg/_0491_ ), .B(\myreg/_2176_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0961_ ) );
MUX2_X1 \myreg/_5298_ ( .A(\myreg/_0502_ ), .B(\myreg/_2178_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0962_ ) );
MUX2_X1 \myreg/_5299_ ( .A(\myreg/_0505_ ), .B(\myreg/_2180_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0963_ ) );
MUX2_X1 \myreg/_5300_ ( .A(\myreg/_0506_ ), .B(\myreg/_2182_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0964_ ) );
MUX2_X1 \myreg/_5301_ ( .A(\myreg/_0507_ ), .B(\myreg/_2184_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0965_ ) );
MUX2_X1 \myreg/_5302_ ( .A(\myreg/_0508_ ), .B(\myreg/_2186_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0966_ ) );
MUX2_X1 \myreg/_5303_ ( .A(\myreg/_0509_ ), .B(\myreg/_2188_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0967_ ) );
MUX2_X1 \myreg/_5304_ ( .A(\myreg/_0510_ ), .B(\myreg/_2190_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0968_ ) );
MUX2_X1 \myreg/_5305_ ( .A(\myreg/_0511_ ), .B(\myreg/_2192_ ), .S(\myreg/_2333_ ), .Z(\myreg/_0969_ ) );
BUF_X4 \myreg/_5306_ ( .A(\myreg/_2332_ ), .Z(\myreg/_2334_ ) );
MUX2_X1 \myreg/_5307_ ( .A(\myreg/_0481_ ), .B(\myreg/_2195_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0970_ ) );
MUX2_X1 \myreg/_5308_ ( .A(\myreg/_0482_ ), .B(\myreg/_2198_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0971_ ) );
MUX2_X1 \myreg/_5309_ ( .A(\myreg/_0483_ ), .B(\myreg/_2200_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0972_ ) );
MUX2_X1 \myreg/_5310_ ( .A(\myreg/_0484_ ), .B(\myreg/_2202_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0973_ ) );
MUX2_X1 \myreg/_5311_ ( .A(\myreg/_0485_ ), .B(\myreg/_2204_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0974_ ) );
MUX2_X1 \myreg/_5312_ ( .A(\myreg/_0486_ ), .B(\myreg/_2206_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0975_ ) );
MUX2_X1 \myreg/_5313_ ( .A(\myreg/_0487_ ), .B(\myreg/_2208_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0976_ ) );
MUX2_X1 \myreg/_5314_ ( .A(\myreg/_0488_ ), .B(\myreg/_2210_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0977_ ) );
MUX2_X1 \myreg/_5315_ ( .A(\myreg/_0489_ ), .B(\myreg/_2212_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0978_ ) );
MUX2_X1 \myreg/_5316_ ( .A(\myreg/_0490_ ), .B(\myreg/_2214_ ), .S(\myreg/_2334_ ), .Z(\myreg/_0979_ ) );
BUF_X4 \myreg/_5317_ ( .A(\myreg/_2332_ ), .Z(\myreg/_2335_ ) );
MUX2_X1 \myreg/_5318_ ( .A(\myreg/_0492_ ), .B(\myreg/_2217_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0980_ ) );
MUX2_X1 \myreg/_5319_ ( .A(\myreg/_0493_ ), .B(\myreg/_2220_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0981_ ) );
MUX2_X1 \myreg/_5320_ ( .A(\myreg/_0494_ ), .B(\myreg/_2222_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0982_ ) );
MUX2_X1 \myreg/_5321_ ( .A(\myreg/_0495_ ), .B(\myreg/_2224_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0983_ ) );
MUX2_X1 \myreg/_5322_ ( .A(\myreg/_0496_ ), .B(\myreg/_2226_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0984_ ) );
MUX2_X1 \myreg/_5323_ ( .A(\myreg/_0497_ ), .B(\myreg/_2228_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0985_ ) );
MUX2_X1 \myreg/_5324_ ( .A(\myreg/_0498_ ), .B(\myreg/_2230_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0986_ ) );
MUX2_X1 \myreg/_5325_ ( .A(\myreg/_0499_ ), .B(\myreg/_2232_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0987_ ) );
MUX2_X1 \myreg/_5326_ ( .A(\myreg/_0500_ ), .B(\myreg/_2234_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0988_ ) );
MUX2_X1 \myreg/_5327_ ( .A(\myreg/_0501_ ), .B(\myreg/_2236_ ), .S(\myreg/_2335_ ), .Z(\myreg/_0989_ ) );
MUX2_X1 \myreg/_5328_ ( .A(\myreg/_0503_ ), .B(\myreg/_2238_ ), .S(\myreg/_2332_ ), .Z(\myreg/_0990_ ) );
MUX2_X1 \myreg/_5329_ ( .A(\myreg/_0504_ ), .B(\myreg/_2240_ ), .S(\myreg/_2332_ ), .Z(\myreg/_0991_ ) );
NOR2_X4 \myreg/_5330_ ( .A1(\myreg/_2173_ ), .A2(\myreg/_2251_ ), .ZN(\myreg/_2336_ ) );
BUF_X4 \myreg/_5331_ ( .A(\myreg/_2336_ ), .Z(\myreg/_2337_ ) );
MUX2_X1 \myreg/_5332_ ( .A(\myreg/_0352_ ), .B(\myreg/_2167_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0992_ ) );
MUX2_X1 \myreg/_5333_ ( .A(\myreg/_0363_ ), .B(\myreg/_2176_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0993_ ) );
MUX2_X1 \myreg/_5334_ ( .A(\myreg/_0374_ ), .B(\myreg/_2178_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0994_ ) );
MUX2_X1 \myreg/_5335_ ( .A(\myreg/_0377_ ), .B(\myreg/_2180_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0995_ ) );
MUX2_X1 \myreg/_5336_ ( .A(\myreg/_0378_ ), .B(\myreg/_2182_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0996_ ) );
MUX2_X1 \myreg/_5337_ ( .A(\myreg/_0379_ ), .B(\myreg/_2184_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0997_ ) );
MUX2_X1 \myreg/_5338_ ( .A(\myreg/_0380_ ), .B(\myreg/_2186_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0998_ ) );
MUX2_X1 \myreg/_5339_ ( .A(\myreg/_0381_ ), .B(\myreg/_2188_ ), .S(\myreg/_2337_ ), .Z(\myreg/_0999_ ) );
MUX2_X1 \myreg/_5340_ ( .A(\myreg/_0382_ ), .B(\myreg/_2190_ ), .S(\myreg/_2337_ ), .Z(\myreg/_1000_ ) );
MUX2_X1 \myreg/_5341_ ( .A(\myreg/_0383_ ), .B(\myreg/_2192_ ), .S(\myreg/_2337_ ), .Z(\myreg/_1001_ ) );
BUF_X4 \myreg/_5342_ ( .A(\myreg/_2336_ ), .Z(\myreg/_2338_ ) );
MUX2_X1 \myreg/_5343_ ( .A(\myreg/_0353_ ), .B(\myreg/_2195_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1002_ ) );
MUX2_X1 \myreg/_5344_ ( .A(\myreg/_0354_ ), .B(\myreg/_2198_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1003_ ) );
MUX2_X1 \myreg/_5345_ ( .A(\myreg/_0355_ ), .B(\myreg/_2200_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1004_ ) );
MUX2_X1 \myreg/_5346_ ( .A(\myreg/_0356_ ), .B(\myreg/_2202_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1005_ ) );
MUX2_X1 \myreg/_5347_ ( .A(\myreg/_0357_ ), .B(\myreg/_2204_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1006_ ) );
MUX2_X1 \myreg/_5348_ ( .A(\myreg/_0358_ ), .B(\myreg/_2206_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1007_ ) );
MUX2_X1 \myreg/_5349_ ( .A(\myreg/_0359_ ), .B(\myreg/_2208_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1008_ ) );
MUX2_X1 \myreg/_5350_ ( .A(\myreg/_0360_ ), .B(\myreg/_2210_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1009_ ) );
MUX2_X1 \myreg/_5351_ ( .A(\myreg/_0361_ ), .B(\myreg/_2212_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1010_ ) );
MUX2_X1 \myreg/_5352_ ( .A(\myreg/_0362_ ), .B(\myreg/_2214_ ), .S(\myreg/_2338_ ), .Z(\myreg/_1011_ ) );
BUF_X4 \myreg/_5353_ ( .A(\myreg/_2336_ ), .Z(\myreg/_2339_ ) );
MUX2_X1 \myreg/_5354_ ( .A(\myreg/_0364_ ), .B(\myreg/_2217_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1012_ ) );
MUX2_X1 \myreg/_5355_ ( .A(\myreg/_0365_ ), .B(\myreg/_2220_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1013_ ) );
MUX2_X1 \myreg/_5356_ ( .A(\myreg/_0366_ ), .B(\myreg/_2222_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1014_ ) );
MUX2_X1 \myreg/_5357_ ( .A(\myreg/_0367_ ), .B(\myreg/_2224_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1015_ ) );
MUX2_X1 \myreg/_5358_ ( .A(\myreg/_0368_ ), .B(\myreg/_2226_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1016_ ) );
MUX2_X1 \myreg/_5359_ ( .A(\myreg/_0369_ ), .B(\myreg/_2228_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1017_ ) );
MUX2_X1 \myreg/_5360_ ( .A(\myreg/_0370_ ), .B(\myreg/_2230_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1018_ ) );
MUX2_X1 \myreg/_5361_ ( .A(\myreg/_0371_ ), .B(\myreg/_2232_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1019_ ) );
MUX2_X1 \myreg/_5362_ ( .A(\myreg/_0372_ ), .B(\myreg/_2234_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1020_ ) );
MUX2_X1 \myreg/_5363_ ( .A(\myreg/_0373_ ), .B(\myreg/_2236_ ), .S(\myreg/_2339_ ), .Z(\myreg/_1021_ ) );
MUX2_X1 \myreg/_5364_ ( .A(\myreg/_0375_ ), .B(\myreg/_2238_ ), .S(\myreg/_2336_ ), .Z(\myreg/_1022_ ) );
MUX2_X1 \myreg/_5365_ ( .A(\myreg/_0376_ ), .B(\myreg/_2240_ ), .S(\myreg/_2336_ ), .Z(\myreg/_1023_ ) );
DFF_X1 \myreg/_5366_ ( .D(\myreg/_2962_ ), .CK(clock ), .Q(\myreg/Reg[7][0] ), .QN(\myreg/_2961_ ) );
DFF_X1 \myreg/_5367_ ( .D(\myreg/_2963_ ), .CK(clock ), .Q(\myreg/Reg[7][1] ), .QN(\myreg/_2960_ ) );
DFF_X1 \myreg/_5368_ ( .D(\myreg/_2964_ ), .CK(clock ), .Q(\myreg/Reg[7][2] ), .QN(\myreg/_2959_ ) );
DFF_X1 \myreg/_5369_ ( .D(\myreg/_2965_ ), .CK(clock ), .Q(\myreg/Reg[7][3] ), .QN(\myreg/_2958_ ) );
DFF_X1 \myreg/_5370_ ( .D(\myreg/_2966_ ), .CK(clock ), .Q(\myreg/Reg[7][4] ), .QN(\myreg/_2957_ ) );
DFF_X1 \myreg/_5371_ ( .D(\myreg/_2967_ ), .CK(clock ), .Q(\myreg/Reg[7][5] ), .QN(\myreg/_2956_ ) );
DFF_X1 \myreg/_5372_ ( .D(\myreg/_2968_ ), .CK(clock ), .Q(\myreg/Reg[7][6] ), .QN(\myreg/_2955_ ) );
DFF_X1 \myreg/_5373_ ( .D(\myreg/_2969_ ), .CK(clock ), .Q(\myreg/Reg[7][7] ), .QN(\myreg/_2954_ ) );
DFF_X1 \myreg/_5374_ ( .D(\myreg/_2970_ ), .CK(clock ), .Q(\myreg/Reg[7][8] ), .QN(\myreg/_2953_ ) );
DFF_X1 \myreg/_5375_ ( .D(\myreg/_2971_ ), .CK(clock ), .Q(\myreg/Reg[7][9] ), .QN(\myreg/_2952_ ) );
DFF_X1 \myreg/_5376_ ( .D(\myreg/_2972_ ), .CK(clock ), .Q(\myreg/Reg[7][10] ), .QN(\myreg/_2951_ ) );
DFF_X1 \myreg/_5377_ ( .D(\myreg/_2973_ ), .CK(clock ), .Q(\myreg/Reg[7][11] ), .QN(\myreg/_2950_ ) );
DFF_X1 \myreg/_5378_ ( .D(\myreg/_2974_ ), .CK(clock ), .Q(\myreg/Reg[7][12] ), .QN(\myreg/_2949_ ) );
DFF_X1 \myreg/_5379_ ( .D(\myreg/_2975_ ), .CK(clock ), .Q(\myreg/Reg[7][13] ), .QN(\myreg/_2948_ ) );
DFF_X1 \myreg/_5380_ ( .D(\myreg/_2976_ ), .CK(clock ), .Q(\myreg/Reg[7][14] ), .QN(\myreg/_2947_ ) );
DFF_X1 \myreg/_5381_ ( .D(\myreg/_2977_ ), .CK(clock ), .Q(\myreg/Reg[7][15] ), .QN(\myreg/_2946_ ) );
DFF_X1 \myreg/_5382_ ( .D(\myreg/_2978_ ), .CK(clock ), .Q(\myreg/Reg[7][16] ), .QN(\myreg/_2945_ ) );
DFF_X1 \myreg/_5383_ ( .D(\myreg/_2979_ ), .CK(clock ), .Q(\myreg/Reg[7][17] ), .QN(\myreg/_2944_ ) );
DFF_X1 \myreg/_5384_ ( .D(\myreg/_2980_ ), .CK(clock ), .Q(\myreg/Reg[7][18] ), .QN(\myreg/_2943_ ) );
DFF_X1 \myreg/_5385_ ( .D(\myreg/_2981_ ), .CK(clock ), .Q(\myreg/Reg[7][19] ), .QN(\myreg/_2942_ ) );
DFF_X1 \myreg/_5386_ ( .D(\myreg/_2982_ ), .CK(clock ), .Q(\myreg/Reg[7][20] ), .QN(\myreg/_2941_ ) );
DFF_X1 \myreg/_5387_ ( .D(\myreg/_2983_ ), .CK(clock ), .Q(\myreg/Reg[7][21] ), .QN(\myreg/_2940_ ) );
DFF_X1 \myreg/_5388_ ( .D(\myreg/_2984_ ), .CK(clock ), .Q(\myreg/Reg[7][22] ), .QN(\myreg/_2939_ ) );
DFF_X1 \myreg/_5389_ ( .D(\myreg/_2985_ ), .CK(clock ), .Q(\myreg/Reg[7][23] ), .QN(\myreg/_2938_ ) );
DFF_X1 \myreg/_5390_ ( .D(\myreg/_2986_ ), .CK(clock ), .Q(\myreg/Reg[7][24] ), .QN(\myreg/_2937_ ) );
DFF_X1 \myreg/_5391_ ( .D(\myreg/_2987_ ), .CK(clock ), .Q(\myreg/Reg[7][25] ), .QN(\myreg/_2936_ ) );
DFF_X1 \myreg/_5392_ ( .D(\myreg/_2988_ ), .CK(clock ), .Q(\myreg/Reg[7][26] ), .QN(\myreg/_2935_ ) );
DFF_X1 \myreg/_5393_ ( .D(\myreg/_2989_ ), .CK(clock ), .Q(\myreg/Reg[7][27] ), .QN(\myreg/_2934_ ) );
DFF_X1 \myreg/_5394_ ( .D(\myreg/_2990_ ), .CK(clock ), .Q(\myreg/Reg[7][28] ), .QN(\myreg/_2933_ ) );
DFF_X1 \myreg/_5395_ ( .D(\myreg/_2991_ ), .CK(clock ), .Q(\myreg/Reg[7][29] ), .QN(\myreg/_2932_ ) );
DFF_X1 \myreg/_5396_ ( .D(\myreg/_2992_ ), .CK(clock ), .Q(\myreg/Reg[7][30] ), .QN(\myreg/_2931_ ) );
DFF_X1 \myreg/_5397_ ( .D(\myreg/_2993_ ), .CK(clock ), .Q(\myreg/Reg[7][31] ), .QN(\myreg/_2930_ ) );
DFF_X1 \myreg/_5398_ ( .D(\myreg/_2994_ ), .CK(clock ), .Q(\myreg/Reg[2][0] ), .QN(\myreg/_2929_ ) );
DFF_X1 \myreg/_5399_ ( .D(\myreg/_2995_ ), .CK(clock ), .Q(\myreg/Reg[2][1] ), .QN(\myreg/_2928_ ) );
DFF_X1 \myreg/_5400_ ( .D(\myreg/_2996_ ), .CK(clock ), .Q(\myreg/Reg[2][2] ), .QN(\myreg/_2927_ ) );
DFF_X1 \myreg/_5401_ ( .D(\myreg/_2997_ ), .CK(clock ), .Q(\myreg/Reg[2][3] ), .QN(\myreg/_2926_ ) );
DFF_X1 \myreg/_5402_ ( .D(\myreg/_2998_ ), .CK(clock ), .Q(\myreg/Reg[2][4] ), .QN(\myreg/_2925_ ) );
DFF_X1 \myreg/_5403_ ( .D(\myreg/_2999_ ), .CK(clock ), .Q(\myreg/Reg[2][5] ), .QN(\myreg/_2924_ ) );
DFF_X1 \myreg/_5404_ ( .D(\myreg/_3000_ ), .CK(clock ), .Q(\myreg/Reg[2][6] ), .QN(\myreg/_2923_ ) );
DFF_X1 \myreg/_5405_ ( .D(\myreg/_3001_ ), .CK(clock ), .Q(\myreg/Reg[2][7] ), .QN(\myreg/_2922_ ) );
DFF_X1 \myreg/_5406_ ( .D(\myreg/_3002_ ), .CK(clock ), .Q(\myreg/Reg[2][8] ), .QN(\myreg/_2921_ ) );
DFF_X1 \myreg/_5407_ ( .D(\myreg/_3003_ ), .CK(clock ), .Q(\myreg/Reg[2][9] ), .QN(\myreg/_2920_ ) );
DFF_X1 \myreg/_5408_ ( .D(\myreg/_3004_ ), .CK(clock ), .Q(\myreg/Reg[2][10] ), .QN(\myreg/_2919_ ) );
DFF_X1 \myreg/_5409_ ( .D(\myreg/_3005_ ), .CK(clock ), .Q(\myreg/Reg[2][11] ), .QN(\myreg/_2918_ ) );
DFF_X1 \myreg/_5410_ ( .D(\myreg/_3006_ ), .CK(clock ), .Q(\myreg/Reg[2][12] ), .QN(\myreg/_2917_ ) );
DFF_X1 \myreg/_5411_ ( .D(\myreg/_3007_ ), .CK(clock ), .Q(\myreg/Reg[2][13] ), .QN(\myreg/_2916_ ) );
DFF_X1 \myreg/_5412_ ( .D(\myreg/_3008_ ), .CK(clock ), .Q(\myreg/Reg[2][14] ), .QN(\myreg/_2915_ ) );
DFF_X1 \myreg/_5413_ ( .D(\myreg/_3009_ ), .CK(clock ), .Q(\myreg/Reg[2][15] ), .QN(\myreg/_2914_ ) );
DFF_X1 \myreg/_5414_ ( .D(\myreg/_3010_ ), .CK(clock ), .Q(\myreg/Reg[2][16] ), .QN(\myreg/_2913_ ) );
DFF_X1 \myreg/_5415_ ( .D(\myreg/_3011_ ), .CK(clock ), .Q(\myreg/Reg[2][17] ), .QN(\myreg/_2912_ ) );
DFF_X1 \myreg/_5416_ ( .D(\myreg/_3012_ ), .CK(clock ), .Q(\myreg/Reg[2][18] ), .QN(\myreg/_2911_ ) );
DFF_X1 \myreg/_5417_ ( .D(\myreg/_3013_ ), .CK(clock ), .Q(\myreg/Reg[2][19] ), .QN(\myreg/_2910_ ) );
DFF_X1 \myreg/_5418_ ( .D(\myreg/_3014_ ), .CK(clock ), .Q(\myreg/Reg[2][20] ), .QN(\myreg/_2909_ ) );
DFF_X1 \myreg/_5419_ ( .D(\myreg/_3015_ ), .CK(clock ), .Q(\myreg/Reg[2][21] ), .QN(\myreg/_2908_ ) );
DFF_X1 \myreg/_5420_ ( .D(\myreg/_3016_ ), .CK(clock ), .Q(\myreg/Reg[2][22] ), .QN(\myreg/_2907_ ) );
DFF_X1 \myreg/_5421_ ( .D(\myreg/_3017_ ), .CK(clock ), .Q(\myreg/Reg[2][23] ), .QN(\myreg/_2906_ ) );
DFF_X1 \myreg/_5422_ ( .D(\myreg/_3018_ ), .CK(clock ), .Q(\myreg/Reg[2][24] ), .QN(\myreg/_2905_ ) );
DFF_X1 \myreg/_5423_ ( .D(\myreg/_3019_ ), .CK(clock ), .Q(\myreg/Reg[2][25] ), .QN(\myreg/_2904_ ) );
DFF_X1 \myreg/_5424_ ( .D(\myreg/_3020_ ), .CK(clock ), .Q(\myreg/Reg[2][26] ), .QN(\myreg/_2903_ ) );
DFF_X1 \myreg/_5425_ ( .D(\myreg/_3021_ ), .CK(clock ), .Q(\myreg/Reg[2][27] ), .QN(\myreg/_2902_ ) );
DFF_X1 \myreg/_5426_ ( .D(\myreg/_3022_ ), .CK(clock ), .Q(\myreg/Reg[2][28] ), .QN(\myreg/_2901_ ) );
DFF_X1 \myreg/_5427_ ( .D(\myreg/_3023_ ), .CK(clock ), .Q(\myreg/Reg[2][29] ), .QN(\myreg/_2900_ ) );
DFF_X1 \myreg/_5428_ ( .D(\myreg/_3024_ ), .CK(clock ), .Q(\myreg/Reg[2][30] ), .QN(\myreg/_2899_ ) );
DFF_X1 \myreg/_5429_ ( .D(\myreg/_3025_ ), .CK(clock ), .Q(\myreg/Reg[2][31] ), .QN(\myreg/_2898_ ) );
DFF_X1 \myreg/_5430_ ( .D(\myreg/_3026_ ), .CK(clock ), .Q(\myreg/Reg[1][0] ), .QN(\myreg/_2897_ ) );
DFF_X1 \myreg/_5431_ ( .D(\myreg/_3027_ ), .CK(clock ), .Q(\myreg/Reg[1][1] ), .QN(\myreg/_2896_ ) );
DFF_X1 \myreg/_5432_ ( .D(\myreg/_3028_ ), .CK(clock ), .Q(\myreg/Reg[1][2] ), .QN(\myreg/_2895_ ) );
DFF_X1 \myreg/_5433_ ( .D(\myreg/_3029_ ), .CK(clock ), .Q(\myreg/Reg[1][3] ), .QN(\myreg/_2894_ ) );
DFF_X1 \myreg/_5434_ ( .D(\myreg/_3030_ ), .CK(clock ), .Q(\myreg/Reg[1][4] ), .QN(\myreg/_2893_ ) );
DFF_X1 \myreg/_5435_ ( .D(\myreg/_3031_ ), .CK(clock ), .Q(\myreg/Reg[1][5] ), .QN(\myreg/_2892_ ) );
DFF_X1 \myreg/_5436_ ( .D(\myreg/_3032_ ), .CK(clock ), .Q(\myreg/Reg[1][6] ), .QN(\myreg/_2891_ ) );
DFF_X1 \myreg/_5437_ ( .D(\myreg/_3033_ ), .CK(clock ), .Q(\myreg/Reg[1][7] ), .QN(\myreg/_2890_ ) );
DFF_X1 \myreg/_5438_ ( .D(\myreg/_3034_ ), .CK(clock ), .Q(\myreg/Reg[1][8] ), .QN(\myreg/_2889_ ) );
DFF_X1 \myreg/_5439_ ( .D(\myreg/_3035_ ), .CK(clock ), .Q(\myreg/Reg[1][9] ), .QN(\myreg/_2888_ ) );
DFF_X1 \myreg/_5440_ ( .D(\myreg/_3036_ ), .CK(clock ), .Q(\myreg/Reg[1][10] ), .QN(\myreg/_2887_ ) );
DFF_X1 \myreg/_5441_ ( .D(\myreg/_3037_ ), .CK(clock ), .Q(\myreg/Reg[1][11] ), .QN(\myreg/_2886_ ) );
DFF_X1 \myreg/_5442_ ( .D(\myreg/_3038_ ), .CK(clock ), .Q(\myreg/Reg[1][12] ), .QN(\myreg/_2885_ ) );
DFF_X1 \myreg/_5443_ ( .D(\myreg/_3039_ ), .CK(clock ), .Q(\myreg/Reg[1][13] ), .QN(\myreg/_2884_ ) );
DFF_X1 \myreg/_5444_ ( .D(\myreg/_3040_ ), .CK(clock ), .Q(\myreg/Reg[1][14] ), .QN(\myreg/_2883_ ) );
DFF_X1 \myreg/_5445_ ( .D(\myreg/_3041_ ), .CK(clock ), .Q(\myreg/Reg[1][15] ), .QN(\myreg/_2882_ ) );
DFF_X1 \myreg/_5446_ ( .D(\myreg/_3042_ ), .CK(clock ), .Q(\myreg/Reg[1][16] ), .QN(\myreg/_2881_ ) );
DFF_X1 \myreg/_5447_ ( .D(\myreg/_3043_ ), .CK(clock ), .Q(\myreg/Reg[1][17] ), .QN(\myreg/_2880_ ) );
DFF_X1 \myreg/_5448_ ( .D(\myreg/_3044_ ), .CK(clock ), .Q(\myreg/Reg[1][18] ), .QN(\myreg/_2879_ ) );
DFF_X1 \myreg/_5449_ ( .D(\myreg/_3045_ ), .CK(clock ), .Q(\myreg/Reg[1][19] ), .QN(\myreg/_2878_ ) );
DFF_X1 \myreg/_5450_ ( .D(\myreg/_3046_ ), .CK(clock ), .Q(\myreg/Reg[1][20] ), .QN(\myreg/_2877_ ) );
DFF_X1 \myreg/_5451_ ( .D(\myreg/_3047_ ), .CK(clock ), .Q(\myreg/Reg[1][21] ), .QN(\myreg/_2876_ ) );
DFF_X1 \myreg/_5452_ ( .D(\myreg/_3048_ ), .CK(clock ), .Q(\myreg/Reg[1][22] ), .QN(\myreg/_2875_ ) );
DFF_X1 \myreg/_5453_ ( .D(\myreg/_3049_ ), .CK(clock ), .Q(\myreg/Reg[1][23] ), .QN(\myreg/_2874_ ) );
DFF_X1 \myreg/_5454_ ( .D(\myreg/_3050_ ), .CK(clock ), .Q(\myreg/Reg[1][24] ), .QN(\myreg/_2873_ ) );
DFF_X1 \myreg/_5455_ ( .D(\myreg/_3051_ ), .CK(clock ), .Q(\myreg/Reg[1][25] ), .QN(\myreg/_2872_ ) );
DFF_X1 \myreg/_5456_ ( .D(\myreg/_3052_ ), .CK(clock ), .Q(\myreg/Reg[1][26] ), .QN(\myreg/_2871_ ) );
DFF_X1 \myreg/_5457_ ( .D(\myreg/_3053_ ), .CK(clock ), .Q(\myreg/Reg[1][27] ), .QN(\myreg/_2870_ ) );
DFF_X1 \myreg/_5458_ ( .D(\myreg/_3054_ ), .CK(clock ), .Q(\myreg/Reg[1][28] ), .QN(\myreg/_2869_ ) );
DFF_X1 \myreg/_5459_ ( .D(\myreg/_3055_ ), .CK(clock ), .Q(\myreg/Reg[1][29] ), .QN(\myreg/_2868_ ) );
DFF_X1 \myreg/_5460_ ( .D(\myreg/_3056_ ), .CK(clock ), .Q(\myreg/Reg[1][30] ), .QN(\myreg/_2867_ ) );
DFF_X1 \myreg/_5461_ ( .D(\myreg/_3057_ ), .CK(clock ), .Q(\myreg/Reg[1][31] ), .QN(\myreg/_2866_ ) );
DFF_X1 \myreg/_5462_ ( .D(\myreg/_3058_ ), .CK(clock ), .Q(\myreg/Reg[4][0] ), .QN(\myreg/_2865_ ) );
DFF_X1 \myreg/_5463_ ( .D(\myreg/_3059_ ), .CK(clock ), .Q(\myreg/Reg[4][1] ), .QN(\myreg/_2864_ ) );
DFF_X1 \myreg/_5464_ ( .D(\myreg/_3060_ ), .CK(clock ), .Q(\myreg/Reg[4][2] ), .QN(\myreg/_2863_ ) );
DFF_X1 \myreg/_5465_ ( .D(\myreg/_3061_ ), .CK(clock ), .Q(\myreg/Reg[4][3] ), .QN(\myreg/_2862_ ) );
DFF_X1 \myreg/_5466_ ( .D(\myreg/_3062_ ), .CK(clock ), .Q(\myreg/Reg[4][4] ), .QN(\myreg/_2861_ ) );
DFF_X1 \myreg/_5467_ ( .D(\myreg/_3063_ ), .CK(clock ), .Q(\myreg/Reg[4][5] ), .QN(\myreg/_2860_ ) );
DFF_X1 \myreg/_5468_ ( .D(\myreg/_3064_ ), .CK(clock ), .Q(\myreg/Reg[4][6] ), .QN(\myreg/_2859_ ) );
DFF_X1 \myreg/_5469_ ( .D(\myreg/_3065_ ), .CK(clock ), .Q(\myreg/Reg[4][7] ), .QN(\myreg/_2858_ ) );
DFF_X1 \myreg/_5470_ ( .D(\myreg/_3066_ ), .CK(clock ), .Q(\myreg/Reg[4][8] ), .QN(\myreg/_2857_ ) );
DFF_X1 \myreg/_5471_ ( .D(\myreg/_3067_ ), .CK(clock ), .Q(\myreg/Reg[4][9] ), .QN(\myreg/_2856_ ) );
DFF_X1 \myreg/_5472_ ( .D(\myreg/_3068_ ), .CK(clock ), .Q(\myreg/Reg[4][10] ), .QN(\myreg/_2855_ ) );
DFF_X1 \myreg/_5473_ ( .D(\myreg/_3069_ ), .CK(clock ), .Q(\myreg/Reg[4][11] ), .QN(\myreg/_2854_ ) );
DFF_X1 \myreg/_5474_ ( .D(\myreg/_3070_ ), .CK(clock ), .Q(\myreg/Reg[4][12] ), .QN(\myreg/_2853_ ) );
DFF_X1 \myreg/_5475_ ( .D(\myreg/_3071_ ), .CK(clock ), .Q(\myreg/Reg[4][13] ), .QN(\myreg/_2852_ ) );
DFF_X1 \myreg/_5476_ ( .D(\myreg/_3072_ ), .CK(clock ), .Q(\myreg/Reg[4][14] ), .QN(\myreg/_2851_ ) );
DFF_X1 \myreg/_5477_ ( .D(\myreg/_3073_ ), .CK(clock ), .Q(\myreg/Reg[4][15] ), .QN(\myreg/_2850_ ) );
DFF_X1 \myreg/_5478_ ( .D(\myreg/_3074_ ), .CK(clock ), .Q(\myreg/Reg[4][16] ), .QN(\myreg/_2849_ ) );
DFF_X1 \myreg/_5479_ ( .D(\myreg/_3075_ ), .CK(clock ), .Q(\myreg/Reg[4][17] ), .QN(\myreg/_2848_ ) );
DFF_X1 \myreg/_5480_ ( .D(\myreg/_3076_ ), .CK(clock ), .Q(\myreg/Reg[4][18] ), .QN(\myreg/_2847_ ) );
DFF_X1 \myreg/_5481_ ( .D(\myreg/_3077_ ), .CK(clock ), .Q(\myreg/Reg[4][19] ), .QN(\myreg/_2846_ ) );
DFF_X1 \myreg/_5482_ ( .D(\myreg/_3078_ ), .CK(clock ), .Q(\myreg/Reg[4][20] ), .QN(\myreg/_2845_ ) );
DFF_X1 \myreg/_5483_ ( .D(\myreg/_3079_ ), .CK(clock ), .Q(\myreg/Reg[4][21] ), .QN(\myreg/_2844_ ) );
DFF_X1 \myreg/_5484_ ( .D(\myreg/_3080_ ), .CK(clock ), .Q(\myreg/Reg[4][22] ), .QN(\myreg/_2843_ ) );
DFF_X1 \myreg/_5485_ ( .D(\myreg/_3081_ ), .CK(clock ), .Q(\myreg/Reg[4][23] ), .QN(\myreg/_2842_ ) );
DFF_X1 \myreg/_5486_ ( .D(\myreg/_3082_ ), .CK(clock ), .Q(\myreg/Reg[4][24] ), .QN(\myreg/_2841_ ) );
DFF_X1 \myreg/_5487_ ( .D(\myreg/_3083_ ), .CK(clock ), .Q(\myreg/Reg[4][25] ), .QN(\myreg/_2840_ ) );
DFF_X1 \myreg/_5488_ ( .D(\myreg/_3084_ ), .CK(clock ), .Q(\myreg/Reg[4][26] ), .QN(\myreg/_2839_ ) );
DFF_X1 \myreg/_5489_ ( .D(\myreg/_3085_ ), .CK(clock ), .Q(\myreg/Reg[4][27] ), .QN(\myreg/_2838_ ) );
DFF_X1 \myreg/_5490_ ( .D(\myreg/_3086_ ), .CK(clock ), .Q(\myreg/Reg[4][28] ), .QN(\myreg/_2837_ ) );
DFF_X1 \myreg/_5491_ ( .D(\myreg/_3087_ ), .CK(clock ), .Q(\myreg/Reg[4][29] ), .QN(\myreg/_2836_ ) );
DFF_X1 \myreg/_5492_ ( .D(\myreg/_3088_ ), .CK(clock ), .Q(\myreg/Reg[4][30] ), .QN(\myreg/_2835_ ) );
DFF_X1 \myreg/_5493_ ( .D(\myreg/_3089_ ), .CK(clock ), .Q(\myreg/Reg[4][31] ), .QN(\myreg/_2834_ ) );
DFF_X1 \myreg/_5494_ ( .D(\myreg/_3090_ ), .CK(clock ), .Q(\myreg/Reg[3][0] ), .QN(\myreg/_2833_ ) );
DFF_X1 \myreg/_5495_ ( .D(\myreg/_3091_ ), .CK(clock ), .Q(\myreg/Reg[3][1] ), .QN(\myreg/_2832_ ) );
DFF_X1 \myreg/_5496_ ( .D(\myreg/_3092_ ), .CK(clock ), .Q(\myreg/Reg[3][2] ), .QN(\myreg/_2831_ ) );
DFF_X1 \myreg/_5497_ ( .D(\myreg/_3093_ ), .CK(clock ), .Q(\myreg/Reg[3][3] ), .QN(\myreg/_2830_ ) );
DFF_X1 \myreg/_5498_ ( .D(\myreg/_3094_ ), .CK(clock ), .Q(\myreg/Reg[3][4] ), .QN(\myreg/_2829_ ) );
DFF_X1 \myreg/_5499_ ( .D(\myreg/_3095_ ), .CK(clock ), .Q(\myreg/Reg[3][5] ), .QN(\myreg/_2828_ ) );
DFF_X1 \myreg/_5500_ ( .D(\myreg/_3096_ ), .CK(clock ), .Q(\myreg/Reg[3][6] ), .QN(\myreg/_2827_ ) );
DFF_X1 \myreg/_5501_ ( .D(\myreg/_3097_ ), .CK(clock ), .Q(\myreg/Reg[3][7] ), .QN(\myreg/_2826_ ) );
DFF_X1 \myreg/_5502_ ( .D(\myreg/_3098_ ), .CK(clock ), .Q(\myreg/Reg[3][8] ), .QN(\myreg/_2825_ ) );
DFF_X1 \myreg/_5503_ ( .D(\myreg/_3099_ ), .CK(clock ), .Q(\myreg/Reg[3][9] ), .QN(\myreg/_2824_ ) );
DFF_X1 \myreg/_5504_ ( .D(\myreg/_3100_ ), .CK(clock ), .Q(\myreg/Reg[3][10] ), .QN(\myreg/_2823_ ) );
DFF_X1 \myreg/_5505_ ( .D(\myreg/_3101_ ), .CK(clock ), .Q(\myreg/Reg[3][11] ), .QN(\myreg/_2822_ ) );
DFF_X1 \myreg/_5506_ ( .D(\myreg/_3102_ ), .CK(clock ), .Q(\myreg/Reg[3][12] ), .QN(\myreg/_2821_ ) );
DFF_X1 \myreg/_5507_ ( .D(\myreg/_3103_ ), .CK(clock ), .Q(\myreg/Reg[3][13] ), .QN(\myreg/_2820_ ) );
DFF_X1 \myreg/_5508_ ( .D(\myreg/_3104_ ), .CK(clock ), .Q(\myreg/Reg[3][14] ), .QN(\myreg/_2819_ ) );
DFF_X1 \myreg/_5509_ ( .D(\myreg/_3105_ ), .CK(clock ), .Q(\myreg/Reg[3][15] ), .QN(\myreg/_2818_ ) );
DFF_X1 \myreg/_5510_ ( .D(\myreg/_3106_ ), .CK(clock ), .Q(\myreg/Reg[3][16] ), .QN(\myreg/_2817_ ) );
DFF_X1 \myreg/_5511_ ( .D(\myreg/_3107_ ), .CK(clock ), .Q(\myreg/Reg[3][17] ), .QN(\myreg/_2816_ ) );
DFF_X1 \myreg/_5512_ ( .D(\myreg/_3108_ ), .CK(clock ), .Q(\myreg/Reg[3][18] ), .QN(\myreg/_2815_ ) );
DFF_X1 \myreg/_5513_ ( .D(\myreg/_3109_ ), .CK(clock ), .Q(\myreg/Reg[3][19] ), .QN(\myreg/_2814_ ) );
DFF_X1 \myreg/_5514_ ( .D(\myreg/_3110_ ), .CK(clock ), .Q(\myreg/Reg[3][20] ), .QN(\myreg/_2813_ ) );
DFF_X1 \myreg/_5515_ ( .D(\myreg/_3111_ ), .CK(clock ), .Q(\myreg/Reg[3][21] ), .QN(\myreg/_2812_ ) );
DFF_X1 \myreg/_5516_ ( .D(\myreg/_3112_ ), .CK(clock ), .Q(\myreg/Reg[3][22] ), .QN(\myreg/_2811_ ) );
DFF_X1 \myreg/_5517_ ( .D(\myreg/_3113_ ), .CK(clock ), .Q(\myreg/Reg[3][23] ), .QN(\myreg/_2810_ ) );
DFF_X1 \myreg/_5518_ ( .D(\myreg/_3114_ ), .CK(clock ), .Q(\myreg/Reg[3][24] ), .QN(\myreg/_2809_ ) );
DFF_X1 \myreg/_5519_ ( .D(\myreg/_3115_ ), .CK(clock ), .Q(\myreg/Reg[3][25] ), .QN(\myreg/_2808_ ) );
DFF_X1 \myreg/_5520_ ( .D(\myreg/_3116_ ), .CK(clock ), .Q(\myreg/Reg[3][26] ), .QN(\myreg/_2807_ ) );
DFF_X1 \myreg/_5521_ ( .D(\myreg/_3117_ ), .CK(clock ), .Q(\myreg/Reg[3][27] ), .QN(\myreg/_2806_ ) );
DFF_X1 \myreg/_5522_ ( .D(\myreg/_3118_ ), .CK(clock ), .Q(\myreg/Reg[3][28] ), .QN(\myreg/_2805_ ) );
DFF_X1 \myreg/_5523_ ( .D(\myreg/_3119_ ), .CK(clock ), .Q(\myreg/Reg[3][29] ), .QN(\myreg/_2804_ ) );
DFF_X1 \myreg/_5524_ ( .D(\myreg/_3120_ ), .CK(clock ), .Q(\myreg/Reg[3][30] ), .QN(\myreg/_2803_ ) );
DFF_X1 \myreg/_5525_ ( .D(\myreg/_3121_ ), .CK(clock ), .Q(\myreg/Reg[3][31] ), .QN(\myreg/_2802_ ) );
DFF_X1 \myreg/_5526_ ( .D(\myreg/_3122_ ), .CK(clock ), .Q(\myreg/Reg[8][0] ), .QN(\myreg/_2801_ ) );
DFF_X1 \myreg/_5527_ ( .D(\myreg/_3123_ ), .CK(clock ), .Q(\myreg/Reg[8][1] ), .QN(\myreg/_2800_ ) );
DFF_X1 \myreg/_5528_ ( .D(\myreg/_3124_ ), .CK(clock ), .Q(\myreg/Reg[8][2] ), .QN(\myreg/_2799_ ) );
DFF_X1 \myreg/_5529_ ( .D(\myreg/_3125_ ), .CK(clock ), .Q(\myreg/Reg[8][3] ), .QN(\myreg/_2798_ ) );
DFF_X1 \myreg/_5530_ ( .D(\myreg/_3126_ ), .CK(clock ), .Q(\myreg/Reg[8][4] ), .QN(\myreg/_2797_ ) );
DFF_X1 \myreg/_5531_ ( .D(\myreg/_3127_ ), .CK(clock ), .Q(\myreg/Reg[8][5] ), .QN(\myreg/_2796_ ) );
DFF_X1 \myreg/_5532_ ( .D(\myreg/_3128_ ), .CK(clock ), .Q(\myreg/Reg[8][6] ), .QN(\myreg/_2795_ ) );
DFF_X1 \myreg/_5533_ ( .D(\myreg/_3129_ ), .CK(clock ), .Q(\myreg/Reg[8][7] ), .QN(\myreg/_2794_ ) );
DFF_X1 \myreg/_5534_ ( .D(\myreg/_3130_ ), .CK(clock ), .Q(\myreg/Reg[8][8] ), .QN(\myreg/_2793_ ) );
DFF_X1 \myreg/_5535_ ( .D(\myreg/_3131_ ), .CK(clock ), .Q(\myreg/Reg[8][9] ), .QN(\myreg/_2792_ ) );
DFF_X1 \myreg/_5536_ ( .D(\myreg/_3132_ ), .CK(clock ), .Q(\myreg/Reg[8][10] ), .QN(\myreg/_2791_ ) );
DFF_X1 \myreg/_5537_ ( .D(\myreg/_3133_ ), .CK(clock ), .Q(\myreg/Reg[8][11] ), .QN(\myreg/_2790_ ) );
DFF_X1 \myreg/_5538_ ( .D(\myreg/_3134_ ), .CK(clock ), .Q(\myreg/Reg[8][12] ), .QN(\myreg/_2789_ ) );
DFF_X1 \myreg/_5539_ ( .D(\myreg/_3135_ ), .CK(clock ), .Q(\myreg/Reg[8][13] ), .QN(\myreg/_2788_ ) );
DFF_X1 \myreg/_5540_ ( .D(\myreg/_3136_ ), .CK(clock ), .Q(\myreg/Reg[8][14] ), .QN(\myreg/_2787_ ) );
DFF_X1 \myreg/_5541_ ( .D(\myreg/_3137_ ), .CK(clock ), .Q(\myreg/Reg[8][15] ), .QN(\myreg/_2786_ ) );
DFF_X1 \myreg/_5542_ ( .D(\myreg/_3138_ ), .CK(clock ), .Q(\myreg/Reg[8][16] ), .QN(\myreg/_2785_ ) );
DFF_X1 \myreg/_5543_ ( .D(\myreg/_3139_ ), .CK(clock ), .Q(\myreg/Reg[8][17] ), .QN(\myreg/_2784_ ) );
DFF_X1 \myreg/_5544_ ( .D(\myreg/_3140_ ), .CK(clock ), .Q(\myreg/Reg[8][18] ), .QN(\myreg/_2783_ ) );
DFF_X1 \myreg/_5545_ ( .D(\myreg/_3141_ ), .CK(clock ), .Q(\myreg/Reg[8][19] ), .QN(\myreg/_2782_ ) );
DFF_X1 \myreg/_5546_ ( .D(\myreg/_3142_ ), .CK(clock ), .Q(\myreg/Reg[8][20] ), .QN(\myreg/_2781_ ) );
DFF_X1 \myreg/_5547_ ( .D(\myreg/_3143_ ), .CK(clock ), .Q(\myreg/Reg[8][21] ), .QN(\myreg/_2780_ ) );
DFF_X1 \myreg/_5548_ ( .D(\myreg/_3144_ ), .CK(clock ), .Q(\myreg/Reg[8][22] ), .QN(\myreg/_2779_ ) );
DFF_X1 \myreg/_5549_ ( .D(\myreg/_3145_ ), .CK(clock ), .Q(\myreg/Reg[8][23] ), .QN(\myreg/_2778_ ) );
DFF_X1 \myreg/_5550_ ( .D(\myreg/_3146_ ), .CK(clock ), .Q(\myreg/Reg[8][24] ), .QN(\myreg/_2777_ ) );
DFF_X1 \myreg/_5551_ ( .D(\myreg/_3147_ ), .CK(clock ), .Q(\myreg/Reg[8][25] ), .QN(\myreg/_2776_ ) );
DFF_X1 \myreg/_5552_ ( .D(\myreg/_3148_ ), .CK(clock ), .Q(\myreg/Reg[8][26] ), .QN(\myreg/_2775_ ) );
DFF_X1 \myreg/_5553_ ( .D(\myreg/_3149_ ), .CK(clock ), .Q(\myreg/Reg[8][27] ), .QN(\myreg/_2774_ ) );
DFF_X1 \myreg/_5554_ ( .D(\myreg/_3150_ ), .CK(clock ), .Q(\myreg/Reg[8][28] ), .QN(\myreg/_2773_ ) );
DFF_X1 \myreg/_5555_ ( .D(\myreg/_3151_ ), .CK(clock ), .Q(\myreg/Reg[8][29] ), .QN(\myreg/_2772_ ) );
DFF_X1 \myreg/_5556_ ( .D(\myreg/_3152_ ), .CK(clock ), .Q(\myreg/Reg[8][30] ), .QN(\myreg/_2771_ ) );
DFF_X1 \myreg/_5557_ ( .D(\myreg/_3153_ ), .CK(clock ), .Q(\myreg/Reg[8][31] ), .QN(\myreg/_2770_ ) );
DFF_X1 \myreg/_5558_ ( .D(\myreg/_3154_ ), .CK(clock ), .Q(\myreg/Reg[0][0] ), .QN(\myreg/_2769_ ) );
DFF_X1 \myreg/_5559_ ( .D(\myreg/_3155_ ), .CK(clock ), .Q(\myreg/Reg[0][1] ), .QN(\myreg/_2768_ ) );
DFF_X1 \myreg/_5560_ ( .D(\myreg/_3156_ ), .CK(clock ), .Q(\myreg/Reg[0][2] ), .QN(\myreg/_2767_ ) );
DFF_X1 \myreg/_5561_ ( .D(\myreg/_3157_ ), .CK(clock ), .Q(\myreg/Reg[0][3] ), .QN(\myreg/_2766_ ) );
DFF_X1 \myreg/_5562_ ( .D(\myreg/_3158_ ), .CK(clock ), .Q(\myreg/Reg[0][4] ), .QN(\myreg/_2765_ ) );
DFF_X1 \myreg/_5563_ ( .D(\myreg/_3159_ ), .CK(clock ), .Q(\myreg/Reg[0][5] ), .QN(\myreg/_2764_ ) );
DFF_X1 \myreg/_5564_ ( .D(\myreg/_3160_ ), .CK(clock ), .Q(\myreg/Reg[0][6] ), .QN(\myreg/_2763_ ) );
DFF_X1 \myreg/_5565_ ( .D(\myreg/_3161_ ), .CK(clock ), .Q(\myreg/Reg[0][7] ), .QN(\myreg/_2762_ ) );
DFF_X1 \myreg/_5566_ ( .D(\myreg/_3162_ ), .CK(clock ), .Q(\myreg/Reg[0][8] ), .QN(\myreg/_2761_ ) );
DFF_X1 \myreg/_5567_ ( .D(\myreg/_3163_ ), .CK(clock ), .Q(\myreg/Reg[0][9] ), .QN(\myreg/_2760_ ) );
DFF_X1 \myreg/_5568_ ( .D(\myreg/_3164_ ), .CK(clock ), .Q(\myreg/Reg[0][10] ), .QN(\myreg/_2759_ ) );
DFF_X1 \myreg/_5569_ ( .D(\myreg/_3165_ ), .CK(clock ), .Q(\myreg/Reg[0][11] ), .QN(\myreg/_2758_ ) );
DFF_X1 \myreg/_5570_ ( .D(\myreg/_3166_ ), .CK(clock ), .Q(\myreg/Reg[0][12] ), .QN(\myreg/_2757_ ) );
DFF_X1 \myreg/_5571_ ( .D(\myreg/_3167_ ), .CK(clock ), .Q(\myreg/Reg[0][13] ), .QN(\myreg/_2756_ ) );
DFF_X1 \myreg/_5572_ ( .D(\myreg/_3168_ ), .CK(clock ), .Q(\myreg/Reg[0][14] ), .QN(\myreg/_2755_ ) );
DFF_X1 \myreg/_5573_ ( .D(\myreg/_3169_ ), .CK(clock ), .Q(\myreg/Reg[0][15] ), .QN(\myreg/_2754_ ) );
DFF_X1 \myreg/_5574_ ( .D(\myreg/_3170_ ), .CK(clock ), .Q(\myreg/Reg[0][16] ), .QN(\myreg/_2753_ ) );
DFF_X1 \myreg/_5575_ ( .D(\myreg/_3171_ ), .CK(clock ), .Q(\myreg/Reg[0][17] ), .QN(\myreg/_2752_ ) );
DFF_X1 \myreg/_5576_ ( .D(\myreg/_3172_ ), .CK(clock ), .Q(\myreg/Reg[0][18] ), .QN(\myreg/_2751_ ) );
DFF_X1 \myreg/_5577_ ( .D(\myreg/_3173_ ), .CK(clock ), .Q(\myreg/Reg[0][19] ), .QN(\myreg/_2750_ ) );
DFF_X1 \myreg/_5578_ ( .D(\myreg/_3174_ ), .CK(clock ), .Q(\myreg/Reg[0][20] ), .QN(\myreg/_2749_ ) );
DFF_X1 \myreg/_5579_ ( .D(\myreg/_3175_ ), .CK(clock ), .Q(\myreg/Reg[0][21] ), .QN(\myreg/_2748_ ) );
DFF_X1 \myreg/_5580_ ( .D(\myreg/_3176_ ), .CK(clock ), .Q(\myreg/Reg[0][22] ), .QN(\myreg/_2747_ ) );
DFF_X1 \myreg/_5581_ ( .D(\myreg/_3177_ ), .CK(clock ), .Q(\myreg/Reg[0][23] ), .QN(\myreg/_2746_ ) );
DFF_X1 \myreg/_5582_ ( .D(\myreg/_3178_ ), .CK(clock ), .Q(\myreg/Reg[0][24] ), .QN(\myreg/_2745_ ) );
DFF_X1 \myreg/_5583_ ( .D(\myreg/_3179_ ), .CK(clock ), .Q(\myreg/Reg[0][25] ), .QN(\myreg/_2744_ ) );
DFF_X1 \myreg/_5584_ ( .D(\myreg/_3180_ ), .CK(clock ), .Q(\myreg/Reg[0][26] ), .QN(\myreg/_2743_ ) );
DFF_X1 \myreg/_5585_ ( .D(\myreg/_3181_ ), .CK(clock ), .Q(\myreg/Reg[0][27] ), .QN(\myreg/_2742_ ) );
DFF_X1 \myreg/_5586_ ( .D(\myreg/_3182_ ), .CK(clock ), .Q(\myreg/Reg[0][28] ), .QN(\myreg/_2741_ ) );
DFF_X1 \myreg/_5587_ ( .D(\myreg/_3183_ ), .CK(clock ), .Q(\myreg/Reg[0][29] ), .QN(\myreg/_2740_ ) );
DFF_X1 \myreg/_5588_ ( .D(\myreg/_3184_ ), .CK(clock ), .Q(\myreg/Reg[0][30] ), .QN(\myreg/_2739_ ) );
DFF_X1 \myreg/_5589_ ( .D(\myreg/_3185_ ), .CK(clock ), .Q(\myreg/Reg[0][31] ), .QN(\myreg/_2738_ ) );
DFF_X1 \myreg/_5590_ ( .D(\myreg/_3186_ ), .CK(clock ), .Q(\myreg/Reg[10][0] ), .QN(\myreg/_2737_ ) );
DFF_X1 \myreg/_5591_ ( .D(\myreg/_3187_ ), .CK(clock ), .Q(\myreg/Reg[10][1] ), .QN(\myreg/_2736_ ) );
DFF_X1 \myreg/_5592_ ( .D(\myreg/_3188_ ), .CK(clock ), .Q(\myreg/Reg[10][2] ), .QN(\myreg/_2735_ ) );
DFF_X1 \myreg/_5593_ ( .D(\myreg/_3189_ ), .CK(clock ), .Q(\myreg/Reg[10][3] ), .QN(\myreg/_2734_ ) );
DFF_X1 \myreg/_5594_ ( .D(\myreg/_3190_ ), .CK(clock ), .Q(\myreg/Reg[10][4] ), .QN(\myreg/_2733_ ) );
DFF_X1 \myreg/_5595_ ( .D(\myreg/_3191_ ), .CK(clock ), .Q(\myreg/Reg[10][5] ), .QN(\myreg/_2732_ ) );
DFF_X1 \myreg/_5596_ ( .D(\myreg/_3192_ ), .CK(clock ), .Q(\myreg/Reg[10][6] ), .QN(\myreg/_2731_ ) );
DFF_X1 \myreg/_5597_ ( .D(\myreg/_3193_ ), .CK(clock ), .Q(\myreg/Reg[10][7] ), .QN(\myreg/_2730_ ) );
DFF_X1 \myreg/_5598_ ( .D(\myreg/_3194_ ), .CK(clock ), .Q(\myreg/Reg[10][8] ), .QN(\myreg/_2729_ ) );
DFF_X1 \myreg/_5599_ ( .D(\myreg/_3195_ ), .CK(clock ), .Q(\myreg/Reg[10][9] ), .QN(\myreg/_2728_ ) );
DFF_X1 \myreg/_5600_ ( .D(\myreg/_3196_ ), .CK(clock ), .Q(\myreg/Reg[10][10] ), .QN(\myreg/_2727_ ) );
DFF_X1 \myreg/_5601_ ( .D(\myreg/_3197_ ), .CK(clock ), .Q(\myreg/Reg[10][11] ), .QN(\myreg/_2726_ ) );
DFF_X1 \myreg/_5602_ ( .D(\myreg/_3198_ ), .CK(clock ), .Q(\myreg/Reg[10][12] ), .QN(\myreg/_2725_ ) );
DFF_X1 \myreg/_5603_ ( .D(\myreg/_3199_ ), .CK(clock ), .Q(\myreg/Reg[10][13] ), .QN(\myreg/_2724_ ) );
DFF_X1 \myreg/_5604_ ( .D(\myreg/_3200_ ), .CK(clock ), .Q(\myreg/Reg[10][14] ), .QN(\myreg/_2723_ ) );
DFF_X1 \myreg/_5605_ ( .D(\myreg/_3201_ ), .CK(clock ), .Q(\myreg/Reg[10][15] ), .QN(\myreg/_2722_ ) );
DFF_X1 \myreg/_5606_ ( .D(\myreg/_3202_ ), .CK(clock ), .Q(\myreg/Reg[10][16] ), .QN(\myreg/_2721_ ) );
DFF_X1 \myreg/_5607_ ( .D(\myreg/_3203_ ), .CK(clock ), .Q(\myreg/Reg[10][17] ), .QN(\myreg/_2720_ ) );
DFF_X1 \myreg/_5608_ ( .D(\myreg/_3204_ ), .CK(clock ), .Q(\myreg/Reg[10][18] ), .QN(\myreg/_2719_ ) );
DFF_X1 \myreg/_5609_ ( .D(\myreg/_3205_ ), .CK(clock ), .Q(\myreg/Reg[10][19] ), .QN(\myreg/_2718_ ) );
DFF_X1 \myreg/_5610_ ( .D(\myreg/_3206_ ), .CK(clock ), .Q(\myreg/Reg[10][20] ), .QN(\myreg/_2717_ ) );
DFF_X1 \myreg/_5611_ ( .D(\myreg/_3207_ ), .CK(clock ), .Q(\myreg/Reg[10][21] ), .QN(\myreg/_2716_ ) );
DFF_X1 \myreg/_5612_ ( .D(\myreg/_3208_ ), .CK(clock ), .Q(\myreg/Reg[10][22] ), .QN(\myreg/_2715_ ) );
DFF_X1 \myreg/_5613_ ( .D(\myreg/_3209_ ), .CK(clock ), .Q(\myreg/Reg[10][23] ), .QN(\myreg/_2714_ ) );
DFF_X1 \myreg/_5614_ ( .D(\myreg/_3210_ ), .CK(clock ), .Q(\myreg/Reg[10][24] ), .QN(\myreg/_2713_ ) );
DFF_X1 \myreg/_5615_ ( .D(\myreg/_3211_ ), .CK(clock ), .Q(\myreg/Reg[10][25] ), .QN(\myreg/_2712_ ) );
DFF_X1 \myreg/_5616_ ( .D(\myreg/_3212_ ), .CK(clock ), .Q(\myreg/Reg[10][26] ), .QN(\myreg/_2711_ ) );
DFF_X1 \myreg/_5617_ ( .D(\myreg/_3213_ ), .CK(clock ), .Q(\myreg/Reg[10][27] ), .QN(\myreg/_2710_ ) );
DFF_X1 \myreg/_5618_ ( .D(\myreg/_3214_ ), .CK(clock ), .Q(\myreg/Reg[10][28] ), .QN(\myreg/_2709_ ) );
DFF_X1 \myreg/_5619_ ( .D(\myreg/_3215_ ), .CK(clock ), .Q(\myreg/Reg[10][29] ), .QN(\myreg/_2708_ ) );
DFF_X1 \myreg/_5620_ ( .D(\myreg/_3216_ ), .CK(clock ), .Q(\myreg/Reg[10][30] ), .QN(\myreg/_2707_ ) );
DFF_X1 \myreg/_5621_ ( .D(\myreg/_3217_ ), .CK(clock ), .Q(\myreg/Reg[10][31] ), .QN(\myreg/_2706_ ) );
DFF_X1 \myreg/_5622_ ( .D(\myreg/_3218_ ), .CK(clock ), .Q(\myreg/Reg[11][0] ), .QN(\myreg/_2705_ ) );
DFF_X1 \myreg/_5623_ ( .D(\myreg/_3219_ ), .CK(clock ), .Q(\myreg/Reg[11][1] ), .QN(\myreg/_2704_ ) );
DFF_X1 \myreg/_5624_ ( .D(\myreg/_3220_ ), .CK(clock ), .Q(\myreg/Reg[11][2] ), .QN(\myreg/_2703_ ) );
DFF_X1 \myreg/_5625_ ( .D(\myreg/_3221_ ), .CK(clock ), .Q(\myreg/Reg[11][3] ), .QN(\myreg/_2702_ ) );
DFF_X1 \myreg/_5626_ ( .D(\myreg/_3222_ ), .CK(clock ), .Q(\myreg/Reg[11][4] ), .QN(\myreg/_2701_ ) );
DFF_X1 \myreg/_5627_ ( .D(\myreg/_3223_ ), .CK(clock ), .Q(\myreg/Reg[11][5] ), .QN(\myreg/_2700_ ) );
DFF_X1 \myreg/_5628_ ( .D(\myreg/_3224_ ), .CK(clock ), .Q(\myreg/Reg[11][6] ), .QN(\myreg/_2699_ ) );
DFF_X1 \myreg/_5629_ ( .D(\myreg/_3225_ ), .CK(clock ), .Q(\myreg/Reg[11][7] ), .QN(\myreg/_2698_ ) );
DFF_X1 \myreg/_5630_ ( .D(\myreg/_3226_ ), .CK(clock ), .Q(\myreg/Reg[11][8] ), .QN(\myreg/_2697_ ) );
DFF_X1 \myreg/_5631_ ( .D(\myreg/_3227_ ), .CK(clock ), .Q(\myreg/Reg[11][9] ), .QN(\myreg/_2696_ ) );
DFF_X1 \myreg/_5632_ ( .D(\myreg/_3228_ ), .CK(clock ), .Q(\myreg/Reg[11][10] ), .QN(\myreg/_2695_ ) );
DFF_X1 \myreg/_5633_ ( .D(\myreg/_3229_ ), .CK(clock ), .Q(\myreg/Reg[11][11] ), .QN(\myreg/_2694_ ) );
DFF_X1 \myreg/_5634_ ( .D(\myreg/_3230_ ), .CK(clock ), .Q(\myreg/Reg[11][12] ), .QN(\myreg/_2693_ ) );
DFF_X1 \myreg/_5635_ ( .D(\myreg/_3231_ ), .CK(clock ), .Q(\myreg/Reg[11][13] ), .QN(\myreg/_2692_ ) );
DFF_X1 \myreg/_5636_ ( .D(\myreg/_3232_ ), .CK(clock ), .Q(\myreg/Reg[11][14] ), .QN(\myreg/_2691_ ) );
DFF_X1 \myreg/_5637_ ( .D(\myreg/_3233_ ), .CK(clock ), .Q(\myreg/Reg[11][15] ), .QN(\myreg/_2690_ ) );
DFF_X1 \myreg/_5638_ ( .D(\myreg/_3234_ ), .CK(clock ), .Q(\myreg/Reg[11][16] ), .QN(\myreg/_2689_ ) );
DFF_X1 \myreg/_5639_ ( .D(\myreg/_3235_ ), .CK(clock ), .Q(\myreg/Reg[11][17] ), .QN(\myreg/_2688_ ) );
DFF_X1 \myreg/_5640_ ( .D(\myreg/_3236_ ), .CK(clock ), .Q(\myreg/Reg[11][18] ), .QN(\myreg/_2687_ ) );
DFF_X1 \myreg/_5641_ ( .D(\myreg/_3237_ ), .CK(clock ), .Q(\myreg/Reg[11][19] ), .QN(\myreg/_2686_ ) );
DFF_X1 \myreg/_5642_ ( .D(\myreg/_3238_ ), .CK(clock ), .Q(\myreg/Reg[11][20] ), .QN(\myreg/_2685_ ) );
DFF_X1 \myreg/_5643_ ( .D(\myreg/_3239_ ), .CK(clock ), .Q(\myreg/Reg[11][21] ), .QN(\myreg/_2684_ ) );
DFF_X1 \myreg/_5644_ ( .D(\myreg/_3240_ ), .CK(clock ), .Q(\myreg/Reg[11][22] ), .QN(\myreg/_2683_ ) );
DFF_X1 \myreg/_5645_ ( .D(\myreg/_3241_ ), .CK(clock ), .Q(\myreg/Reg[11][23] ), .QN(\myreg/_2682_ ) );
DFF_X1 \myreg/_5646_ ( .D(\myreg/_3242_ ), .CK(clock ), .Q(\myreg/Reg[11][24] ), .QN(\myreg/_2681_ ) );
DFF_X1 \myreg/_5647_ ( .D(\myreg/_3243_ ), .CK(clock ), .Q(\myreg/Reg[11][25] ), .QN(\myreg/_2680_ ) );
DFF_X1 \myreg/_5648_ ( .D(\myreg/_3244_ ), .CK(clock ), .Q(\myreg/Reg[11][26] ), .QN(\myreg/_2679_ ) );
DFF_X1 \myreg/_5649_ ( .D(\myreg/_3245_ ), .CK(clock ), .Q(\myreg/Reg[11][27] ), .QN(\myreg/_2678_ ) );
DFF_X1 \myreg/_5650_ ( .D(\myreg/_3246_ ), .CK(clock ), .Q(\myreg/Reg[11][28] ), .QN(\myreg/_2677_ ) );
DFF_X1 \myreg/_5651_ ( .D(\myreg/_3247_ ), .CK(clock ), .Q(\myreg/Reg[11][29] ), .QN(\myreg/_2676_ ) );
DFF_X1 \myreg/_5652_ ( .D(\myreg/_3248_ ), .CK(clock ), .Q(\myreg/Reg[11][30] ), .QN(\myreg/_2675_ ) );
DFF_X1 \myreg/_5653_ ( .D(\myreg/_3249_ ), .CK(clock ), .Q(\myreg/Reg[11][31] ), .QN(\myreg/_2674_ ) );
DFF_X1 \myreg/_5654_ ( .D(\myreg/_3250_ ), .CK(clock ), .Q(\myreg/Reg[12][0] ), .QN(\myreg/_2673_ ) );
DFF_X1 \myreg/_5655_ ( .D(\myreg/_3251_ ), .CK(clock ), .Q(\myreg/Reg[12][1] ), .QN(\myreg/_2672_ ) );
DFF_X1 \myreg/_5656_ ( .D(\myreg/_3252_ ), .CK(clock ), .Q(\myreg/Reg[12][2] ), .QN(\myreg/_2671_ ) );
DFF_X1 \myreg/_5657_ ( .D(\myreg/_3253_ ), .CK(clock ), .Q(\myreg/Reg[12][3] ), .QN(\myreg/_2670_ ) );
DFF_X1 \myreg/_5658_ ( .D(\myreg/_3254_ ), .CK(clock ), .Q(\myreg/Reg[12][4] ), .QN(\myreg/_2669_ ) );
DFF_X1 \myreg/_5659_ ( .D(\myreg/_3255_ ), .CK(clock ), .Q(\myreg/Reg[12][5] ), .QN(\myreg/_2668_ ) );
DFF_X1 \myreg/_5660_ ( .D(\myreg/_3256_ ), .CK(clock ), .Q(\myreg/Reg[12][6] ), .QN(\myreg/_2667_ ) );
DFF_X1 \myreg/_5661_ ( .D(\myreg/_3257_ ), .CK(clock ), .Q(\myreg/Reg[12][7] ), .QN(\myreg/_2666_ ) );
DFF_X1 \myreg/_5662_ ( .D(\myreg/_3258_ ), .CK(clock ), .Q(\myreg/Reg[12][8] ), .QN(\myreg/_2665_ ) );
DFF_X1 \myreg/_5663_ ( .D(\myreg/_3259_ ), .CK(clock ), .Q(\myreg/Reg[12][9] ), .QN(\myreg/_2664_ ) );
DFF_X1 \myreg/_5664_ ( .D(\myreg/_3260_ ), .CK(clock ), .Q(\myreg/Reg[12][10] ), .QN(\myreg/_2663_ ) );
DFF_X1 \myreg/_5665_ ( .D(\myreg/_3261_ ), .CK(clock ), .Q(\myreg/Reg[12][11] ), .QN(\myreg/_2662_ ) );
DFF_X1 \myreg/_5666_ ( .D(\myreg/_3262_ ), .CK(clock ), .Q(\myreg/Reg[12][12] ), .QN(\myreg/_2661_ ) );
DFF_X1 \myreg/_5667_ ( .D(\myreg/_3263_ ), .CK(clock ), .Q(\myreg/Reg[12][13] ), .QN(\myreg/_2660_ ) );
DFF_X1 \myreg/_5668_ ( .D(\myreg/_3264_ ), .CK(clock ), .Q(\myreg/Reg[12][14] ), .QN(\myreg/_2659_ ) );
DFF_X1 \myreg/_5669_ ( .D(\myreg/_3265_ ), .CK(clock ), .Q(\myreg/Reg[12][15] ), .QN(\myreg/_2658_ ) );
DFF_X1 \myreg/_5670_ ( .D(\myreg/_3266_ ), .CK(clock ), .Q(\myreg/Reg[12][16] ), .QN(\myreg/_2657_ ) );
DFF_X1 \myreg/_5671_ ( .D(\myreg/_3267_ ), .CK(clock ), .Q(\myreg/Reg[12][17] ), .QN(\myreg/_2656_ ) );
DFF_X1 \myreg/_5672_ ( .D(\myreg/_3268_ ), .CK(clock ), .Q(\myreg/Reg[12][18] ), .QN(\myreg/_2655_ ) );
DFF_X1 \myreg/_5673_ ( .D(\myreg/_3269_ ), .CK(clock ), .Q(\myreg/Reg[12][19] ), .QN(\myreg/_2654_ ) );
DFF_X1 \myreg/_5674_ ( .D(\myreg/_3270_ ), .CK(clock ), .Q(\myreg/Reg[12][20] ), .QN(\myreg/_2653_ ) );
DFF_X1 \myreg/_5675_ ( .D(\myreg/_3271_ ), .CK(clock ), .Q(\myreg/Reg[12][21] ), .QN(\myreg/_2652_ ) );
DFF_X1 \myreg/_5676_ ( .D(\myreg/_3272_ ), .CK(clock ), .Q(\myreg/Reg[12][22] ), .QN(\myreg/_2651_ ) );
DFF_X1 \myreg/_5677_ ( .D(\myreg/_3273_ ), .CK(clock ), .Q(\myreg/Reg[12][23] ), .QN(\myreg/_2650_ ) );
DFF_X1 \myreg/_5678_ ( .D(\myreg/_3274_ ), .CK(clock ), .Q(\myreg/Reg[12][24] ), .QN(\myreg/_2649_ ) );
DFF_X1 \myreg/_5679_ ( .D(\myreg/_3275_ ), .CK(clock ), .Q(\myreg/Reg[12][25] ), .QN(\myreg/_2648_ ) );
DFF_X1 \myreg/_5680_ ( .D(\myreg/_3276_ ), .CK(clock ), .Q(\myreg/Reg[12][26] ), .QN(\myreg/_2647_ ) );
DFF_X1 \myreg/_5681_ ( .D(\myreg/_3277_ ), .CK(clock ), .Q(\myreg/Reg[12][27] ), .QN(\myreg/_2646_ ) );
DFF_X1 \myreg/_5682_ ( .D(\myreg/_3278_ ), .CK(clock ), .Q(\myreg/Reg[12][28] ), .QN(\myreg/_2645_ ) );
DFF_X1 \myreg/_5683_ ( .D(\myreg/_3279_ ), .CK(clock ), .Q(\myreg/Reg[12][29] ), .QN(\myreg/_2644_ ) );
DFF_X1 \myreg/_5684_ ( .D(\myreg/_3280_ ), .CK(clock ), .Q(\myreg/Reg[12][30] ), .QN(\myreg/_2643_ ) );
DFF_X1 \myreg/_5685_ ( .D(\myreg/_3281_ ), .CK(clock ), .Q(\myreg/Reg[12][31] ), .QN(\myreg/_2642_ ) );
DFF_X1 \myreg/_5686_ ( .D(\myreg/_3282_ ), .CK(clock ), .Q(\myreg/Reg[13][0] ), .QN(\myreg/_2641_ ) );
DFF_X1 \myreg/_5687_ ( .D(\myreg/_3283_ ), .CK(clock ), .Q(\myreg/Reg[13][1] ), .QN(\myreg/_2640_ ) );
DFF_X1 \myreg/_5688_ ( .D(\myreg/_3284_ ), .CK(clock ), .Q(\myreg/Reg[13][2] ), .QN(\myreg/_2639_ ) );
DFF_X1 \myreg/_5689_ ( .D(\myreg/_3285_ ), .CK(clock ), .Q(\myreg/Reg[13][3] ), .QN(\myreg/_2638_ ) );
DFF_X1 \myreg/_5690_ ( .D(\myreg/_3286_ ), .CK(clock ), .Q(\myreg/Reg[13][4] ), .QN(\myreg/_2637_ ) );
DFF_X1 \myreg/_5691_ ( .D(\myreg/_3287_ ), .CK(clock ), .Q(\myreg/Reg[13][5] ), .QN(\myreg/_2636_ ) );
DFF_X1 \myreg/_5692_ ( .D(\myreg/_3288_ ), .CK(clock ), .Q(\myreg/Reg[13][6] ), .QN(\myreg/_2635_ ) );
DFF_X1 \myreg/_5693_ ( .D(\myreg/_3289_ ), .CK(clock ), .Q(\myreg/Reg[13][7] ), .QN(\myreg/_2634_ ) );
DFF_X1 \myreg/_5694_ ( .D(\myreg/_3290_ ), .CK(clock ), .Q(\myreg/Reg[13][8] ), .QN(\myreg/_2633_ ) );
DFF_X1 \myreg/_5695_ ( .D(\myreg/_3291_ ), .CK(clock ), .Q(\myreg/Reg[13][9] ), .QN(\myreg/_2632_ ) );
DFF_X1 \myreg/_5696_ ( .D(\myreg/_3292_ ), .CK(clock ), .Q(\myreg/Reg[13][10] ), .QN(\myreg/_2631_ ) );
DFF_X1 \myreg/_5697_ ( .D(\myreg/_3293_ ), .CK(clock ), .Q(\myreg/Reg[13][11] ), .QN(\myreg/_2630_ ) );
DFF_X1 \myreg/_5698_ ( .D(\myreg/_3294_ ), .CK(clock ), .Q(\myreg/Reg[13][12] ), .QN(\myreg/_2629_ ) );
DFF_X1 \myreg/_5699_ ( .D(\myreg/_3295_ ), .CK(clock ), .Q(\myreg/Reg[13][13] ), .QN(\myreg/_2628_ ) );
DFF_X1 \myreg/_5700_ ( .D(\myreg/_3296_ ), .CK(clock ), .Q(\myreg/Reg[13][14] ), .QN(\myreg/_2627_ ) );
DFF_X1 \myreg/_5701_ ( .D(\myreg/_3297_ ), .CK(clock ), .Q(\myreg/Reg[13][15] ), .QN(\myreg/_2626_ ) );
DFF_X1 \myreg/_5702_ ( .D(\myreg/_3298_ ), .CK(clock ), .Q(\myreg/Reg[13][16] ), .QN(\myreg/_2625_ ) );
DFF_X1 \myreg/_5703_ ( .D(\myreg/_3299_ ), .CK(clock ), .Q(\myreg/Reg[13][17] ), .QN(\myreg/_2624_ ) );
DFF_X1 \myreg/_5704_ ( .D(\myreg/_3300_ ), .CK(clock ), .Q(\myreg/Reg[13][18] ), .QN(\myreg/_2623_ ) );
DFF_X1 \myreg/_5705_ ( .D(\myreg/_3301_ ), .CK(clock ), .Q(\myreg/Reg[13][19] ), .QN(\myreg/_2622_ ) );
DFF_X1 \myreg/_5706_ ( .D(\myreg/_3302_ ), .CK(clock ), .Q(\myreg/Reg[13][20] ), .QN(\myreg/_2621_ ) );
DFF_X1 \myreg/_5707_ ( .D(\myreg/_3303_ ), .CK(clock ), .Q(\myreg/Reg[13][21] ), .QN(\myreg/_2620_ ) );
DFF_X1 \myreg/_5708_ ( .D(\myreg/_3304_ ), .CK(clock ), .Q(\myreg/Reg[13][22] ), .QN(\myreg/_2619_ ) );
DFF_X1 \myreg/_5709_ ( .D(\myreg/_3305_ ), .CK(clock ), .Q(\myreg/Reg[13][23] ), .QN(\myreg/_2618_ ) );
DFF_X1 \myreg/_5710_ ( .D(\myreg/_3306_ ), .CK(clock ), .Q(\myreg/Reg[13][24] ), .QN(\myreg/_2617_ ) );
DFF_X1 \myreg/_5711_ ( .D(\myreg/_3307_ ), .CK(clock ), .Q(\myreg/Reg[13][25] ), .QN(\myreg/_2616_ ) );
DFF_X1 \myreg/_5712_ ( .D(\myreg/_3308_ ), .CK(clock ), .Q(\myreg/Reg[13][26] ), .QN(\myreg/_2615_ ) );
DFF_X1 \myreg/_5713_ ( .D(\myreg/_3309_ ), .CK(clock ), .Q(\myreg/Reg[13][27] ), .QN(\myreg/_2614_ ) );
DFF_X1 \myreg/_5714_ ( .D(\myreg/_3310_ ), .CK(clock ), .Q(\myreg/Reg[13][28] ), .QN(\myreg/_2613_ ) );
DFF_X1 \myreg/_5715_ ( .D(\myreg/_3311_ ), .CK(clock ), .Q(\myreg/Reg[13][29] ), .QN(\myreg/_2612_ ) );
DFF_X1 \myreg/_5716_ ( .D(\myreg/_3312_ ), .CK(clock ), .Q(\myreg/Reg[13][30] ), .QN(\myreg/_2611_ ) );
DFF_X1 \myreg/_5717_ ( .D(\myreg/_3313_ ), .CK(clock ), .Q(\myreg/Reg[13][31] ), .QN(\myreg/_2610_ ) );
DFF_X1 \myreg/_5718_ ( .D(\myreg/_3314_ ), .CK(clock ), .Q(\myreg/Reg[14][0] ), .QN(\myreg/_2609_ ) );
DFF_X1 \myreg/_5719_ ( .D(\myreg/_3315_ ), .CK(clock ), .Q(\myreg/Reg[14][1] ), .QN(\myreg/_2608_ ) );
DFF_X1 \myreg/_5720_ ( .D(\myreg/_3316_ ), .CK(clock ), .Q(\myreg/Reg[14][2] ), .QN(\myreg/_2607_ ) );
DFF_X1 \myreg/_5721_ ( .D(\myreg/_3317_ ), .CK(clock ), .Q(\myreg/Reg[14][3] ), .QN(\myreg/_2606_ ) );
DFF_X1 \myreg/_5722_ ( .D(\myreg/_3318_ ), .CK(clock ), .Q(\myreg/Reg[14][4] ), .QN(\myreg/_2605_ ) );
DFF_X1 \myreg/_5723_ ( .D(\myreg/_3319_ ), .CK(clock ), .Q(\myreg/Reg[14][5] ), .QN(\myreg/_2604_ ) );
DFF_X1 \myreg/_5724_ ( .D(\myreg/_3320_ ), .CK(clock ), .Q(\myreg/Reg[14][6] ), .QN(\myreg/_2603_ ) );
DFF_X1 \myreg/_5725_ ( .D(\myreg/_3321_ ), .CK(clock ), .Q(\myreg/Reg[14][7] ), .QN(\myreg/_2602_ ) );
DFF_X1 \myreg/_5726_ ( .D(\myreg/_3322_ ), .CK(clock ), .Q(\myreg/Reg[14][8] ), .QN(\myreg/_2601_ ) );
DFF_X1 \myreg/_5727_ ( .D(\myreg/_3323_ ), .CK(clock ), .Q(\myreg/Reg[14][9] ), .QN(\myreg/_2600_ ) );
DFF_X1 \myreg/_5728_ ( .D(\myreg/_3324_ ), .CK(clock ), .Q(\myreg/Reg[14][10] ), .QN(\myreg/_2599_ ) );
DFF_X1 \myreg/_5729_ ( .D(\myreg/_3325_ ), .CK(clock ), .Q(\myreg/Reg[14][11] ), .QN(\myreg/_2598_ ) );
DFF_X1 \myreg/_5730_ ( .D(\myreg/_3326_ ), .CK(clock ), .Q(\myreg/Reg[14][12] ), .QN(\myreg/_2597_ ) );
DFF_X1 \myreg/_5731_ ( .D(\myreg/_3327_ ), .CK(clock ), .Q(\myreg/Reg[14][13] ), .QN(\myreg/_2596_ ) );
DFF_X1 \myreg/_5732_ ( .D(\myreg/_3328_ ), .CK(clock ), .Q(\myreg/Reg[14][14] ), .QN(\myreg/_2595_ ) );
DFF_X1 \myreg/_5733_ ( .D(\myreg/_3329_ ), .CK(clock ), .Q(\myreg/Reg[14][15] ), .QN(\myreg/_2594_ ) );
DFF_X1 \myreg/_5734_ ( .D(\myreg/_3330_ ), .CK(clock ), .Q(\myreg/Reg[14][16] ), .QN(\myreg/_2593_ ) );
DFF_X1 \myreg/_5735_ ( .D(\myreg/_3331_ ), .CK(clock ), .Q(\myreg/Reg[14][17] ), .QN(\myreg/_2592_ ) );
DFF_X1 \myreg/_5736_ ( .D(\myreg/_3332_ ), .CK(clock ), .Q(\myreg/Reg[14][18] ), .QN(\myreg/_2591_ ) );
DFF_X1 \myreg/_5737_ ( .D(\myreg/_3333_ ), .CK(clock ), .Q(\myreg/Reg[14][19] ), .QN(\myreg/_2590_ ) );
DFF_X1 \myreg/_5738_ ( .D(\myreg/_3334_ ), .CK(clock ), .Q(\myreg/Reg[14][20] ), .QN(\myreg/_2589_ ) );
DFF_X1 \myreg/_5739_ ( .D(\myreg/_3335_ ), .CK(clock ), .Q(\myreg/Reg[14][21] ), .QN(\myreg/_2588_ ) );
DFF_X1 \myreg/_5740_ ( .D(\myreg/_3336_ ), .CK(clock ), .Q(\myreg/Reg[14][22] ), .QN(\myreg/_2587_ ) );
DFF_X1 \myreg/_5741_ ( .D(\myreg/_3337_ ), .CK(clock ), .Q(\myreg/Reg[14][23] ), .QN(\myreg/_2586_ ) );
DFF_X1 \myreg/_5742_ ( .D(\myreg/_3338_ ), .CK(clock ), .Q(\myreg/Reg[14][24] ), .QN(\myreg/_2585_ ) );
DFF_X1 \myreg/_5743_ ( .D(\myreg/_3339_ ), .CK(clock ), .Q(\myreg/Reg[14][25] ), .QN(\myreg/_2584_ ) );
DFF_X1 \myreg/_5744_ ( .D(\myreg/_3340_ ), .CK(clock ), .Q(\myreg/Reg[14][26] ), .QN(\myreg/_2583_ ) );
DFF_X1 \myreg/_5745_ ( .D(\myreg/_3341_ ), .CK(clock ), .Q(\myreg/Reg[14][27] ), .QN(\myreg/_2582_ ) );
DFF_X1 \myreg/_5746_ ( .D(\myreg/_3342_ ), .CK(clock ), .Q(\myreg/Reg[14][28] ), .QN(\myreg/_2581_ ) );
DFF_X1 \myreg/_5747_ ( .D(\myreg/_3343_ ), .CK(clock ), .Q(\myreg/Reg[14][29] ), .QN(\myreg/_2580_ ) );
DFF_X1 \myreg/_5748_ ( .D(\myreg/_3344_ ), .CK(clock ), .Q(\myreg/Reg[14][30] ), .QN(\myreg/_2579_ ) );
DFF_X1 \myreg/_5749_ ( .D(\myreg/_3345_ ), .CK(clock ), .Q(\myreg/Reg[14][31] ), .QN(\myreg/_2578_ ) );
DFF_X1 \myreg/_5750_ ( .D(\myreg/_3346_ ), .CK(clock ), .Q(\myreg/Reg[6][0] ), .QN(\myreg/_2577_ ) );
DFF_X1 \myreg/_5751_ ( .D(\myreg/_3347_ ), .CK(clock ), .Q(\myreg/Reg[6][1] ), .QN(\myreg/_2576_ ) );
DFF_X1 \myreg/_5752_ ( .D(\myreg/_3348_ ), .CK(clock ), .Q(\myreg/Reg[6][2] ), .QN(\myreg/_2575_ ) );
DFF_X1 \myreg/_5753_ ( .D(\myreg/_3349_ ), .CK(clock ), .Q(\myreg/Reg[6][3] ), .QN(\myreg/_2574_ ) );
DFF_X1 \myreg/_5754_ ( .D(\myreg/_3350_ ), .CK(clock ), .Q(\myreg/Reg[6][4] ), .QN(\myreg/_2573_ ) );
DFF_X1 \myreg/_5755_ ( .D(\myreg/_3351_ ), .CK(clock ), .Q(\myreg/Reg[6][5] ), .QN(\myreg/_2572_ ) );
DFF_X1 \myreg/_5756_ ( .D(\myreg/_3352_ ), .CK(clock ), .Q(\myreg/Reg[6][6] ), .QN(\myreg/_2571_ ) );
DFF_X1 \myreg/_5757_ ( .D(\myreg/_3353_ ), .CK(clock ), .Q(\myreg/Reg[6][7] ), .QN(\myreg/_2570_ ) );
DFF_X1 \myreg/_5758_ ( .D(\myreg/_3354_ ), .CK(clock ), .Q(\myreg/Reg[6][8] ), .QN(\myreg/_2569_ ) );
DFF_X1 \myreg/_5759_ ( .D(\myreg/_3355_ ), .CK(clock ), .Q(\myreg/Reg[6][9] ), .QN(\myreg/_2568_ ) );
DFF_X1 \myreg/_5760_ ( .D(\myreg/_3356_ ), .CK(clock ), .Q(\myreg/Reg[6][10] ), .QN(\myreg/_2567_ ) );
DFF_X1 \myreg/_5761_ ( .D(\myreg/_3357_ ), .CK(clock ), .Q(\myreg/Reg[6][11] ), .QN(\myreg/_2566_ ) );
DFF_X1 \myreg/_5762_ ( .D(\myreg/_3358_ ), .CK(clock ), .Q(\myreg/Reg[6][12] ), .QN(\myreg/_2565_ ) );
DFF_X1 \myreg/_5763_ ( .D(\myreg/_3359_ ), .CK(clock ), .Q(\myreg/Reg[6][13] ), .QN(\myreg/_2564_ ) );
DFF_X1 \myreg/_5764_ ( .D(\myreg/_3360_ ), .CK(clock ), .Q(\myreg/Reg[6][14] ), .QN(\myreg/_2563_ ) );
DFF_X1 \myreg/_5765_ ( .D(\myreg/_3361_ ), .CK(clock ), .Q(\myreg/Reg[6][15] ), .QN(\myreg/_2562_ ) );
DFF_X1 \myreg/_5766_ ( .D(\myreg/_3362_ ), .CK(clock ), .Q(\myreg/Reg[6][16] ), .QN(\myreg/_2561_ ) );
DFF_X1 \myreg/_5767_ ( .D(\myreg/_3363_ ), .CK(clock ), .Q(\myreg/Reg[6][17] ), .QN(\myreg/_2560_ ) );
DFF_X1 \myreg/_5768_ ( .D(\myreg/_3364_ ), .CK(clock ), .Q(\myreg/Reg[6][18] ), .QN(\myreg/_2559_ ) );
DFF_X1 \myreg/_5769_ ( .D(\myreg/_3365_ ), .CK(clock ), .Q(\myreg/Reg[6][19] ), .QN(\myreg/_2558_ ) );
DFF_X1 \myreg/_5770_ ( .D(\myreg/_3366_ ), .CK(clock ), .Q(\myreg/Reg[6][20] ), .QN(\myreg/_2557_ ) );
DFF_X1 \myreg/_5771_ ( .D(\myreg/_3367_ ), .CK(clock ), .Q(\myreg/Reg[6][21] ), .QN(\myreg/_2556_ ) );
DFF_X1 \myreg/_5772_ ( .D(\myreg/_3368_ ), .CK(clock ), .Q(\myreg/Reg[6][22] ), .QN(\myreg/_2555_ ) );
DFF_X1 \myreg/_5773_ ( .D(\myreg/_3369_ ), .CK(clock ), .Q(\myreg/Reg[6][23] ), .QN(\myreg/_2554_ ) );
DFF_X1 \myreg/_5774_ ( .D(\myreg/_3370_ ), .CK(clock ), .Q(\myreg/Reg[6][24] ), .QN(\myreg/_2553_ ) );
DFF_X1 \myreg/_5775_ ( .D(\myreg/_3371_ ), .CK(clock ), .Q(\myreg/Reg[6][25] ), .QN(\myreg/_2552_ ) );
DFF_X1 \myreg/_5776_ ( .D(\myreg/_3372_ ), .CK(clock ), .Q(\myreg/Reg[6][26] ), .QN(\myreg/_2551_ ) );
DFF_X1 \myreg/_5777_ ( .D(\myreg/_3373_ ), .CK(clock ), .Q(\myreg/Reg[6][27] ), .QN(\myreg/_2550_ ) );
DFF_X1 \myreg/_5778_ ( .D(\myreg/_3374_ ), .CK(clock ), .Q(\myreg/Reg[6][28] ), .QN(\myreg/_2549_ ) );
DFF_X1 \myreg/_5779_ ( .D(\myreg/_3375_ ), .CK(clock ), .Q(\myreg/Reg[6][29] ), .QN(\myreg/_2548_ ) );
DFF_X1 \myreg/_5780_ ( .D(\myreg/_3376_ ), .CK(clock ), .Q(\myreg/Reg[6][30] ), .QN(\myreg/_2547_ ) );
DFF_X1 \myreg/_5781_ ( .D(\myreg/_3377_ ), .CK(clock ), .Q(\myreg/Reg[6][31] ), .QN(\myreg/_2546_ ) );
DFF_X1 \myreg/_5782_ ( .D(\myreg/_3378_ ), .CK(clock ), .Q(\myreg/Reg[15][0] ), .QN(\myreg/_2545_ ) );
DFF_X1 \myreg/_5783_ ( .D(\myreg/_3379_ ), .CK(clock ), .Q(\myreg/Reg[15][1] ), .QN(\myreg/_2544_ ) );
DFF_X1 \myreg/_5784_ ( .D(\myreg/_3380_ ), .CK(clock ), .Q(\myreg/Reg[15][2] ), .QN(\myreg/_2543_ ) );
DFF_X1 \myreg/_5785_ ( .D(\myreg/_3381_ ), .CK(clock ), .Q(\myreg/Reg[15][3] ), .QN(\myreg/_2542_ ) );
DFF_X1 \myreg/_5786_ ( .D(\myreg/_3382_ ), .CK(clock ), .Q(\myreg/Reg[15][4] ), .QN(\myreg/_2541_ ) );
DFF_X1 \myreg/_5787_ ( .D(\myreg/_3383_ ), .CK(clock ), .Q(\myreg/Reg[15][5] ), .QN(\myreg/_2540_ ) );
DFF_X1 \myreg/_5788_ ( .D(\myreg/_3384_ ), .CK(clock ), .Q(\myreg/Reg[15][6] ), .QN(\myreg/_2539_ ) );
DFF_X1 \myreg/_5789_ ( .D(\myreg/_3385_ ), .CK(clock ), .Q(\myreg/Reg[15][7] ), .QN(\myreg/_2538_ ) );
DFF_X1 \myreg/_5790_ ( .D(\myreg/_3386_ ), .CK(clock ), .Q(\myreg/Reg[15][8] ), .QN(\myreg/_2537_ ) );
DFF_X1 \myreg/_5791_ ( .D(\myreg/_3387_ ), .CK(clock ), .Q(\myreg/Reg[15][9] ), .QN(\myreg/_2536_ ) );
DFF_X1 \myreg/_5792_ ( .D(\myreg/_3388_ ), .CK(clock ), .Q(\myreg/Reg[15][10] ), .QN(\myreg/_2535_ ) );
DFF_X1 \myreg/_5793_ ( .D(\myreg/_3389_ ), .CK(clock ), .Q(\myreg/Reg[15][11] ), .QN(\myreg/_2534_ ) );
DFF_X1 \myreg/_5794_ ( .D(\myreg/_3390_ ), .CK(clock ), .Q(\myreg/Reg[15][12] ), .QN(\myreg/_2533_ ) );
DFF_X1 \myreg/_5795_ ( .D(\myreg/_3391_ ), .CK(clock ), .Q(\myreg/Reg[15][13] ), .QN(\myreg/_2532_ ) );
DFF_X1 \myreg/_5796_ ( .D(\myreg/_3392_ ), .CK(clock ), .Q(\myreg/Reg[15][14] ), .QN(\myreg/_2531_ ) );
DFF_X1 \myreg/_5797_ ( .D(\myreg/_3393_ ), .CK(clock ), .Q(\myreg/Reg[15][15] ), .QN(\myreg/_2530_ ) );
DFF_X1 \myreg/_5798_ ( .D(\myreg/_3394_ ), .CK(clock ), .Q(\myreg/Reg[15][16] ), .QN(\myreg/_2529_ ) );
DFF_X1 \myreg/_5799_ ( .D(\myreg/_3395_ ), .CK(clock ), .Q(\myreg/Reg[15][17] ), .QN(\myreg/_2528_ ) );
DFF_X1 \myreg/_5800_ ( .D(\myreg/_3396_ ), .CK(clock ), .Q(\myreg/Reg[15][18] ), .QN(\myreg/_2527_ ) );
DFF_X1 \myreg/_5801_ ( .D(\myreg/_3397_ ), .CK(clock ), .Q(\myreg/Reg[15][19] ), .QN(\myreg/_2526_ ) );
DFF_X1 \myreg/_5802_ ( .D(\myreg/_3398_ ), .CK(clock ), .Q(\myreg/Reg[15][20] ), .QN(\myreg/_2525_ ) );
DFF_X1 \myreg/_5803_ ( .D(\myreg/_3399_ ), .CK(clock ), .Q(\myreg/Reg[15][21] ), .QN(\myreg/_2524_ ) );
DFF_X1 \myreg/_5804_ ( .D(\myreg/_3400_ ), .CK(clock ), .Q(\myreg/Reg[15][22] ), .QN(\myreg/_2523_ ) );
DFF_X1 \myreg/_5805_ ( .D(\myreg/_3401_ ), .CK(clock ), .Q(\myreg/Reg[15][23] ), .QN(\myreg/_2522_ ) );
DFF_X1 \myreg/_5806_ ( .D(\myreg/_3402_ ), .CK(clock ), .Q(\myreg/Reg[15][24] ), .QN(\myreg/_2521_ ) );
DFF_X1 \myreg/_5807_ ( .D(\myreg/_3403_ ), .CK(clock ), .Q(\myreg/Reg[15][25] ), .QN(\myreg/_2520_ ) );
DFF_X1 \myreg/_5808_ ( .D(\myreg/_3404_ ), .CK(clock ), .Q(\myreg/Reg[15][26] ), .QN(\myreg/_2519_ ) );
DFF_X1 \myreg/_5809_ ( .D(\myreg/_3405_ ), .CK(clock ), .Q(\myreg/Reg[15][27] ), .QN(\myreg/_2518_ ) );
DFF_X1 \myreg/_5810_ ( .D(\myreg/_3406_ ), .CK(clock ), .Q(\myreg/Reg[15][28] ), .QN(\myreg/_2517_ ) );
DFF_X1 \myreg/_5811_ ( .D(\myreg/_3407_ ), .CK(clock ), .Q(\myreg/Reg[15][29] ), .QN(\myreg/_2516_ ) );
DFF_X1 \myreg/_5812_ ( .D(\myreg/_3408_ ), .CK(clock ), .Q(\myreg/Reg[15][30] ), .QN(\myreg/_2515_ ) );
DFF_X1 \myreg/_5813_ ( .D(\myreg/_3409_ ), .CK(clock ), .Q(\myreg/Reg[15][31] ), .QN(\myreg/_2514_ ) );
DFF_X1 \myreg/_5814_ ( .D(\myreg/_3410_ ), .CK(clock ), .Q(\myreg/Reg[9][0] ), .QN(\myreg/_2513_ ) );
DFF_X1 \myreg/_5815_ ( .D(\myreg/_3411_ ), .CK(clock ), .Q(\myreg/Reg[9][1] ), .QN(\myreg/_2512_ ) );
DFF_X1 \myreg/_5816_ ( .D(\myreg/_3412_ ), .CK(clock ), .Q(\myreg/Reg[9][2] ), .QN(\myreg/_2511_ ) );
DFF_X1 \myreg/_5817_ ( .D(\myreg/_3413_ ), .CK(clock ), .Q(\myreg/Reg[9][3] ), .QN(\myreg/_2510_ ) );
DFF_X1 \myreg/_5818_ ( .D(\myreg/_3414_ ), .CK(clock ), .Q(\myreg/Reg[9][4] ), .QN(\myreg/_2509_ ) );
DFF_X1 \myreg/_5819_ ( .D(\myreg/_3415_ ), .CK(clock ), .Q(\myreg/Reg[9][5] ), .QN(\myreg/_2508_ ) );
DFF_X1 \myreg/_5820_ ( .D(\myreg/_3416_ ), .CK(clock ), .Q(\myreg/Reg[9][6] ), .QN(\myreg/_2507_ ) );
DFF_X1 \myreg/_5821_ ( .D(\myreg/_3417_ ), .CK(clock ), .Q(\myreg/Reg[9][7] ), .QN(\myreg/_2506_ ) );
DFF_X1 \myreg/_5822_ ( .D(\myreg/_3418_ ), .CK(clock ), .Q(\myreg/Reg[9][8] ), .QN(\myreg/_2505_ ) );
DFF_X1 \myreg/_5823_ ( .D(\myreg/_3419_ ), .CK(clock ), .Q(\myreg/Reg[9][9] ), .QN(\myreg/_2504_ ) );
DFF_X1 \myreg/_5824_ ( .D(\myreg/_3420_ ), .CK(clock ), .Q(\myreg/Reg[9][10] ), .QN(\myreg/_2503_ ) );
DFF_X1 \myreg/_5825_ ( .D(\myreg/_3421_ ), .CK(clock ), .Q(\myreg/Reg[9][11] ), .QN(\myreg/_2502_ ) );
DFF_X1 \myreg/_5826_ ( .D(\myreg/_3422_ ), .CK(clock ), .Q(\myreg/Reg[9][12] ), .QN(\myreg/_2501_ ) );
DFF_X1 \myreg/_5827_ ( .D(\myreg/_3423_ ), .CK(clock ), .Q(\myreg/Reg[9][13] ), .QN(\myreg/_2500_ ) );
DFF_X1 \myreg/_5828_ ( .D(\myreg/_3424_ ), .CK(clock ), .Q(\myreg/Reg[9][14] ), .QN(\myreg/_2499_ ) );
DFF_X1 \myreg/_5829_ ( .D(\myreg/_3425_ ), .CK(clock ), .Q(\myreg/Reg[9][15] ), .QN(\myreg/_2498_ ) );
DFF_X1 \myreg/_5830_ ( .D(\myreg/_3426_ ), .CK(clock ), .Q(\myreg/Reg[9][16] ), .QN(\myreg/_2497_ ) );
DFF_X1 \myreg/_5831_ ( .D(\myreg/_3427_ ), .CK(clock ), .Q(\myreg/Reg[9][17] ), .QN(\myreg/_2496_ ) );
DFF_X1 \myreg/_5832_ ( .D(\myreg/_3428_ ), .CK(clock ), .Q(\myreg/Reg[9][18] ), .QN(\myreg/_2495_ ) );
DFF_X1 \myreg/_5833_ ( .D(\myreg/_3429_ ), .CK(clock ), .Q(\myreg/Reg[9][19] ), .QN(\myreg/_2494_ ) );
DFF_X1 \myreg/_5834_ ( .D(\myreg/_3430_ ), .CK(clock ), .Q(\myreg/Reg[9][20] ), .QN(\myreg/_2493_ ) );
DFF_X1 \myreg/_5835_ ( .D(\myreg/_3431_ ), .CK(clock ), .Q(\myreg/Reg[9][21] ), .QN(\myreg/_2492_ ) );
DFF_X1 \myreg/_5836_ ( .D(\myreg/_3432_ ), .CK(clock ), .Q(\myreg/Reg[9][22] ), .QN(\myreg/_2491_ ) );
DFF_X1 \myreg/_5837_ ( .D(\myreg/_3433_ ), .CK(clock ), .Q(\myreg/Reg[9][23] ), .QN(\myreg/_2490_ ) );
DFF_X1 \myreg/_5838_ ( .D(\myreg/_3434_ ), .CK(clock ), .Q(\myreg/Reg[9][24] ), .QN(\myreg/_2489_ ) );
DFF_X1 \myreg/_5839_ ( .D(\myreg/_3435_ ), .CK(clock ), .Q(\myreg/Reg[9][25] ), .QN(\myreg/_2488_ ) );
DFF_X1 \myreg/_5840_ ( .D(\myreg/_3436_ ), .CK(clock ), .Q(\myreg/Reg[9][26] ), .QN(\myreg/_2487_ ) );
DFF_X1 \myreg/_5841_ ( .D(\myreg/_3437_ ), .CK(clock ), .Q(\myreg/Reg[9][27] ), .QN(\myreg/_2486_ ) );
DFF_X1 \myreg/_5842_ ( .D(\myreg/_3438_ ), .CK(clock ), .Q(\myreg/Reg[9][28] ), .QN(\myreg/_2485_ ) );
DFF_X1 \myreg/_5843_ ( .D(\myreg/_3439_ ), .CK(clock ), .Q(\myreg/Reg[9][29] ), .QN(\myreg/_2484_ ) );
DFF_X1 \myreg/_5844_ ( .D(\myreg/_3440_ ), .CK(clock ), .Q(\myreg/Reg[9][30] ), .QN(\myreg/_2483_ ) );
DFF_X1 \myreg/_5845_ ( .D(\myreg/_3441_ ), .CK(clock ), .Q(\myreg/Reg[9][31] ), .QN(\myreg/_2482_ ) );
DFF_X1 \myreg/_5846_ ( .D(\myreg/_3442_ ), .CK(clock ), .Q(\myreg/Reg[5][0] ), .QN(\myreg/_2481_ ) );
DFF_X1 \myreg/_5847_ ( .D(\myreg/_3443_ ), .CK(clock ), .Q(\myreg/Reg[5][1] ), .QN(\myreg/_2480_ ) );
DFF_X1 \myreg/_5848_ ( .D(\myreg/_3444_ ), .CK(clock ), .Q(\myreg/Reg[5][2] ), .QN(\myreg/_2479_ ) );
DFF_X1 \myreg/_5849_ ( .D(\myreg/_3445_ ), .CK(clock ), .Q(\myreg/Reg[5][3] ), .QN(\myreg/_2478_ ) );
DFF_X1 \myreg/_5850_ ( .D(\myreg/_3446_ ), .CK(clock ), .Q(\myreg/Reg[5][4] ), .QN(\myreg/_2477_ ) );
DFF_X1 \myreg/_5851_ ( .D(\myreg/_3447_ ), .CK(clock ), .Q(\myreg/Reg[5][5] ), .QN(\myreg/_2476_ ) );
DFF_X1 \myreg/_5852_ ( .D(\myreg/_3448_ ), .CK(clock ), .Q(\myreg/Reg[5][6] ), .QN(\myreg/_2475_ ) );
DFF_X1 \myreg/_5853_ ( .D(\myreg/_3449_ ), .CK(clock ), .Q(\myreg/Reg[5][7] ), .QN(\myreg/_2474_ ) );
DFF_X1 \myreg/_5854_ ( .D(\myreg/_3450_ ), .CK(clock ), .Q(\myreg/Reg[5][8] ), .QN(\myreg/_2473_ ) );
DFF_X1 \myreg/_5855_ ( .D(\myreg/_3451_ ), .CK(clock ), .Q(\myreg/Reg[5][9] ), .QN(\myreg/_2472_ ) );
DFF_X1 \myreg/_5856_ ( .D(\myreg/_3452_ ), .CK(clock ), .Q(\myreg/Reg[5][10] ), .QN(\myreg/_2471_ ) );
DFF_X1 \myreg/_5857_ ( .D(\myreg/_3453_ ), .CK(clock ), .Q(\myreg/Reg[5][11] ), .QN(\myreg/_2470_ ) );
DFF_X1 \myreg/_5858_ ( .D(\myreg/_3454_ ), .CK(clock ), .Q(\myreg/Reg[5][12] ), .QN(\myreg/_2469_ ) );
DFF_X1 \myreg/_5859_ ( .D(\myreg/_3455_ ), .CK(clock ), .Q(\myreg/Reg[5][13] ), .QN(\myreg/_2468_ ) );
DFF_X1 \myreg/_5860_ ( .D(\myreg/_3456_ ), .CK(clock ), .Q(\myreg/Reg[5][14] ), .QN(\myreg/_2467_ ) );
DFF_X1 \myreg/_5861_ ( .D(\myreg/_3457_ ), .CK(clock ), .Q(\myreg/Reg[5][15] ), .QN(\myreg/_2466_ ) );
DFF_X1 \myreg/_5862_ ( .D(\myreg/_3458_ ), .CK(clock ), .Q(\myreg/Reg[5][16] ), .QN(\myreg/_2465_ ) );
DFF_X1 \myreg/_5863_ ( .D(\myreg/_3459_ ), .CK(clock ), .Q(\myreg/Reg[5][17] ), .QN(\myreg/_2464_ ) );
DFF_X1 \myreg/_5864_ ( .D(\myreg/_3460_ ), .CK(clock ), .Q(\myreg/Reg[5][18] ), .QN(\myreg/_2463_ ) );
DFF_X1 \myreg/_5865_ ( .D(\myreg/_3461_ ), .CK(clock ), .Q(\myreg/Reg[5][19] ), .QN(\myreg/_2462_ ) );
DFF_X1 \myreg/_5866_ ( .D(\myreg/_3462_ ), .CK(clock ), .Q(\myreg/Reg[5][20] ), .QN(\myreg/_2461_ ) );
DFF_X1 \myreg/_5867_ ( .D(\myreg/_3463_ ), .CK(clock ), .Q(\myreg/Reg[5][21] ), .QN(\myreg/_2460_ ) );
DFF_X1 \myreg/_5868_ ( .D(\myreg/_3464_ ), .CK(clock ), .Q(\myreg/Reg[5][22] ), .QN(\myreg/_2459_ ) );
DFF_X1 \myreg/_5869_ ( .D(\myreg/_3465_ ), .CK(clock ), .Q(\myreg/Reg[5][23] ), .QN(\myreg/_2458_ ) );
DFF_X1 \myreg/_5870_ ( .D(\myreg/_3466_ ), .CK(clock ), .Q(\myreg/Reg[5][24] ), .QN(\myreg/_2457_ ) );
DFF_X1 \myreg/_5871_ ( .D(\myreg/_3467_ ), .CK(clock ), .Q(\myreg/Reg[5][25] ), .QN(\myreg/_2456_ ) );
DFF_X1 \myreg/_5872_ ( .D(\myreg/_3468_ ), .CK(clock ), .Q(\myreg/Reg[5][26] ), .QN(\myreg/_2455_ ) );
DFF_X1 \myreg/_5873_ ( .D(\myreg/_3469_ ), .CK(clock ), .Q(\myreg/Reg[5][27] ), .QN(\myreg/_2454_ ) );
DFF_X1 \myreg/_5874_ ( .D(\myreg/_3470_ ), .CK(clock ), .Q(\myreg/Reg[5][28] ), .QN(\myreg/_2453_ ) );
DFF_X1 \myreg/_5875_ ( .D(\myreg/_3471_ ), .CK(clock ), .Q(\myreg/Reg[5][29] ), .QN(\myreg/_2452_ ) );
DFF_X1 \myreg/_5876_ ( .D(\myreg/_3472_ ), .CK(clock ), .Q(\myreg/Reg[5][30] ), .QN(\myreg/_2451_ ) );
DFF_X1 \myreg/_5877_ ( .D(\myreg/_3473_ ), .CK(clock ), .Q(\myreg/Reg[5][31] ), .QN(\myreg/_2450_ ) );
BUF_X1 \myreg/_5878_ ( .A(\LS_WB_waddr_reg [1] ), .Z(\myreg/_2414_ ) );
BUF_X1 \myreg/_5879_ ( .A(\LS_WB_waddr_reg [0] ), .Z(\myreg/_2413_ ) );
BUF_X1 \myreg/_5880_ ( .A(\LS_WB_waddr_reg [3] ), .Z(\myreg/_2416_ ) );
BUF_X1 \myreg/_5881_ ( .A(\LS_WB_waddr_reg [2] ), .Z(\myreg/_2415_ ) );
BUF_X1 \myreg/_5882_ ( .A(LS_WB_wen_reg ), .Z(\myreg/_2449_ ) );
BUF_X1 \myreg/_5883_ ( .A(reset ), .Z(\myreg/_2412_ ) );
BUF_X1 \myreg/_5884_ ( .A(\LS_WB_wdata_reg [0] ), .Z(\myreg/_2417_ ) );
BUF_X1 \myreg/_5885_ ( .A(\LS_WB_wdata_reg [1] ), .Z(\myreg/_2428_ ) );
BUF_X1 \myreg/_5886_ ( .A(\LS_WB_wdata_reg [2] ), .Z(\myreg/_2439_ ) );
BUF_X1 \myreg/_5887_ ( .A(\LS_WB_wdata_reg [3] ), .Z(\myreg/_2442_ ) );
BUF_X1 \myreg/_5888_ ( .A(\LS_WB_wdata_reg [4] ), .Z(\myreg/_2443_ ) );
BUF_X1 \myreg/_5889_ ( .A(\LS_WB_wdata_reg [5] ), .Z(\myreg/_2444_ ) );
BUF_X1 \myreg/_5890_ ( .A(\LS_WB_wdata_reg [6] ), .Z(\myreg/_2445_ ) );
BUF_X1 \myreg/_5891_ ( .A(\LS_WB_wdata_reg [7] ), .Z(\myreg/_2446_ ) );
BUF_X1 \myreg/_5892_ ( .A(\LS_WB_wdata_reg [8] ), .Z(\myreg/_2447_ ) );
BUF_X1 \myreg/_5893_ ( .A(\LS_WB_wdata_reg [9] ), .Z(\myreg/_2448_ ) );
BUF_X1 \myreg/_5894_ ( .A(\LS_WB_wdata_reg [10] ), .Z(\myreg/_2418_ ) );
BUF_X1 \myreg/_5895_ ( .A(\LS_WB_wdata_reg [11] ), .Z(\myreg/_2419_ ) );
BUF_X1 \myreg/_5896_ ( .A(\LS_WB_wdata_reg [12] ), .Z(\myreg/_2420_ ) );
BUF_X1 \myreg/_5897_ ( .A(\LS_WB_wdata_reg [13] ), .Z(\myreg/_2421_ ) );
BUF_X1 \myreg/_5898_ ( .A(\LS_WB_wdata_reg [14] ), .Z(\myreg/_2422_ ) );
BUF_X1 \myreg/_5899_ ( .A(\LS_WB_wdata_reg [15] ), .Z(\myreg/_2423_ ) );
BUF_X1 \myreg/_5900_ ( .A(\LS_WB_wdata_reg [16] ), .Z(\myreg/_2424_ ) );
BUF_X1 \myreg/_5901_ ( .A(\LS_WB_wdata_reg [17] ), .Z(\myreg/_2425_ ) );
BUF_X1 \myreg/_5902_ ( .A(\LS_WB_wdata_reg [18] ), .Z(\myreg/_2426_ ) );
BUF_X1 \myreg/_5903_ ( .A(\LS_WB_wdata_reg [19] ), .Z(\myreg/_2427_ ) );
BUF_X1 \myreg/_5904_ ( .A(\LS_WB_wdata_reg [20] ), .Z(\myreg/_2429_ ) );
BUF_X1 \myreg/_5905_ ( .A(\LS_WB_wdata_reg [21] ), .Z(\myreg/_2430_ ) );
BUF_X1 \myreg/_5906_ ( .A(\LS_WB_wdata_reg [22] ), .Z(\myreg/_2431_ ) );
BUF_X1 \myreg/_5907_ ( .A(\LS_WB_wdata_reg [23] ), .Z(\myreg/_2432_ ) );
BUF_X1 \myreg/_5908_ ( .A(\LS_WB_wdata_reg [24] ), .Z(\myreg/_2433_ ) );
BUF_X1 \myreg/_5909_ ( .A(\LS_WB_wdata_reg [25] ), .Z(\myreg/_2434_ ) );
BUF_X1 \myreg/_5910_ ( .A(\LS_WB_wdata_reg [26] ), .Z(\myreg/_2435_ ) );
BUF_X1 \myreg/_5911_ ( .A(\LS_WB_wdata_reg [27] ), .Z(\myreg/_2436_ ) );
BUF_X1 \myreg/_5912_ ( .A(\LS_WB_wdata_reg [28] ), .Z(\myreg/_2437_ ) );
BUF_X1 \myreg/_5913_ ( .A(\LS_WB_wdata_reg [29] ), .Z(\myreg/_2438_ ) );
BUF_X1 \myreg/_5914_ ( .A(\LS_WB_wdata_reg [30] ), .Z(\myreg/_2440_ ) );
BUF_X1 \myreg/_5915_ ( .A(\LS_WB_wdata_reg [31] ), .Z(\myreg/_2441_ ) );
BUF_X1 \myreg/_5916_ ( .A(\myreg/Reg[0][0] ), .Z(\myreg/_0000_ ) );
BUF_X1 \myreg/_5917_ ( .A(\myreg/Reg[1][0] ), .Z(\myreg/_0224_ ) );
BUF_X1 \myreg/_5918_ ( .A(\ID_EX_rs1 [0] ), .Z(\myreg/_2340_ ) );
BUF_X1 \myreg/_5919_ ( .A(\myreg/Reg[2][0] ), .Z(\myreg/_0256_ ) );
BUF_X1 \myreg/_5920_ ( .A(\myreg/Reg[3][0] ), .Z(\myreg/_0288_ ) );
BUF_X1 \myreg/_5921_ ( .A(\ID_EX_rs1 [1] ), .Z(\myreg/_2341_ ) );
BUF_X1 \myreg/_5922_ ( .A(\myreg/Reg[4][0] ), .Z(\myreg/_0320_ ) );
BUF_X1 \myreg/_5923_ ( .A(\myreg/Reg[5][0] ), .Z(\myreg/_0352_ ) );
BUF_X1 \myreg/_5924_ ( .A(\myreg/Reg[6][0] ), .Z(\myreg/_0384_ ) );
BUF_X1 \myreg/_5925_ ( .A(\myreg/Reg[7][0] ), .Z(\myreg/_0416_ ) );
BUF_X1 \myreg/_5926_ ( .A(\ID_EX_rs1 [2] ), .Z(\myreg/_2342_ ) );
BUF_X1 \myreg/_5927_ ( .A(\myreg/Reg[8][0] ), .Z(\myreg/_0448_ ) );
BUF_X1 \myreg/_5928_ ( .A(\myreg/Reg[9][0] ), .Z(\myreg/_0480_ ) );
BUF_X1 \myreg/_5929_ ( .A(\myreg/Reg[10][0] ), .Z(\myreg/_0032_ ) );
BUF_X1 \myreg/_5930_ ( .A(\myreg/Reg[11][0] ), .Z(\myreg/_0064_ ) );
BUF_X1 \myreg/_5931_ ( .A(\myreg/Reg[12][0] ), .Z(\myreg/_0096_ ) );
BUF_X1 \myreg/_5932_ ( .A(\myreg/Reg[13][0] ), .Z(\myreg/_0128_ ) );
BUF_X1 \myreg/_5933_ ( .A(\myreg/Reg[14][0] ), .Z(\myreg/_0160_ ) );
BUF_X1 \myreg/_5934_ ( .A(\myreg/Reg[15][0] ), .Z(\myreg/_0192_ ) );
BUF_X1 \myreg/_5935_ ( .A(\ID_EX_rs1 [3] ), .Z(\myreg/_2343_ ) );
BUF_X1 \myreg/_5936_ ( .A(\myreg/_2348_ ), .Z(\src1_raw [0] ) );
BUF_X1 \myreg/_5937_ ( .A(\myreg/Reg[0][1] ), .Z(\myreg/_0011_ ) );
BUF_X1 \myreg/_5938_ ( .A(\myreg/Reg[1][1] ), .Z(\myreg/_0235_ ) );
BUF_X1 \myreg/_5939_ ( .A(\myreg/Reg[2][1] ), .Z(\myreg/_0267_ ) );
BUF_X1 \myreg/_5940_ ( .A(\myreg/Reg[3][1] ), .Z(\myreg/_0299_ ) );
BUF_X1 \myreg/_5941_ ( .A(\myreg/Reg[4][1] ), .Z(\myreg/_0331_ ) );
BUF_X1 \myreg/_5942_ ( .A(\myreg/Reg[5][1] ), .Z(\myreg/_0363_ ) );
BUF_X1 \myreg/_5943_ ( .A(\myreg/Reg[6][1] ), .Z(\myreg/_0395_ ) );
BUF_X1 \myreg/_5944_ ( .A(\myreg/Reg[7][1] ), .Z(\myreg/_0427_ ) );
BUF_X1 \myreg/_5945_ ( .A(\myreg/Reg[8][1] ), .Z(\myreg/_0459_ ) );
BUF_X1 \myreg/_5946_ ( .A(\myreg/Reg[9][1] ), .Z(\myreg/_0491_ ) );
BUF_X1 \myreg/_5947_ ( .A(\myreg/Reg[10][1] ), .Z(\myreg/_0043_ ) );
BUF_X1 \myreg/_5948_ ( .A(\myreg/Reg[11][1] ), .Z(\myreg/_0075_ ) );
BUF_X1 \myreg/_5949_ ( .A(\myreg/Reg[12][1] ), .Z(\myreg/_0107_ ) );
BUF_X1 \myreg/_5950_ ( .A(\myreg/Reg[13][1] ), .Z(\myreg/_0139_ ) );
BUF_X1 \myreg/_5951_ ( .A(\myreg/Reg[14][1] ), .Z(\myreg/_0171_ ) );
BUF_X1 \myreg/_5952_ ( .A(\myreg/Reg[15][1] ), .Z(\myreg/_0203_ ) );
BUF_X1 \myreg/_5953_ ( .A(\myreg/_2359_ ), .Z(\src1_raw [1] ) );
BUF_X1 \myreg/_5954_ ( .A(\myreg/Reg[0][2] ), .Z(\myreg/_0022_ ) );
BUF_X1 \myreg/_5955_ ( .A(\myreg/Reg[1][2] ), .Z(\myreg/_0246_ ) );
BUF_X1 \myreg/_5956_ ( .A(\myreg/Reg[2][2] ), .Z(\myreg/_0278_ ) );
BUF_X1 \myreg/_5957_ ( .A(\myreg/Reg[3][2] ), .Z(\myreg/_0310_ ) );
BUF_X1 \myreg/_5958_ ( .A(\myreg/Reg[4][2] ), .Z(\myreg/_0342_ ) );
BUF_X1 \myreg/_5959_ ( .A(\myreg/Reg[5][2] ), .Z(\myreg/_0374_ ) );
BUF_X1 \myreg/_5960_ ( .A(\myreg/Reg[6][2] ), .Z(\myreg/_0406_ ) );
BUF_X1 \myreg/_5961_ ( .A(\myreg/Reg[7][2] ), .Z(\myreg/_0438_ ) );
BUF_X1 \myreg/_5962_ ( .A(\myreg/Reg[8][2] ), .Z(\myreg/_0470_ ) );
BUF_X1 \myreg/_5963_ ( .A(\myreg/Reg[9][2] ), .Z(\myreg/_0502_ ) );
BUF_X1 \myreg/_5964_ ( .A(\myreg/Reg[10][2] ), .Z(\myreg/_0054_ ) );
BUF_X1 \myreg/_5965_ ( .A(\myreg/Reg[11][2] ), .Z(\myreg/_0086_ ) );
BUF_X1 \myreg/_5966_ ( .A(\myreg/Reg[12][2] ), .Z(\myreg/_0118_ ) );
BUF_X1 \myreg/_5967_ ( .A(\myreg/Reg[13][2] ), .Z(\myreg/_0150_ ) );
BUF_X1 \myreg/_5968_ ( .A(\myreg/Reg[14][2] ), .Z(\myreg/_0182_ ) );
BUF_X1 \myreg/_5969_ ( .A(\myreg/Reg[15][2] ), .Z(\myreg/_0214_ ) );
BUF_X1 \myreg/_5970_ ( .A(\myreg/_2370_ ), .Z(\src1_raw [2] ) );
BUF_X1 \myreg/_5971_ ( .A(\myreg/Reg[0][3] ), .Z(\myreg/_0025_ ) );
BUF_X1 \myreg/_5972_ ( .A(\myreg/Reg[1][3] ), .Z(\myreg/_0249_ ) );
BUF_X1 \myreg/_5973_ ( .A(\myreg/Reg[2][3] ), .Z(\myreg/_0281_ ) );
BUF_X1 \myreg/_5974_ ( .A(\myreg/Reg[3][3] ), .Z(\myreg/_0313_ ) );
BUF_X1 \myreg/_5975_ ( .A(\myreg/Reg[4][3] ), .Z(\myreg/_0345_ ) );
BUF_X1 \myreg/_5976_ ( .A(\myreg/Reg[5][3] ), .Z(\myreg/_0377_ ) );
BUF_X1 \myreg/_5977_ ( .A(\myreg/Reg[6][3] ), .Z(\myreg/_0409_ ) );
BUF_X1 \myreg/_5978_ ( .A(\myreg/Reg[7][3] ), .Z(\myreg/_0441_ ) );
BUF_X1 \myreg/_5979_ ( .A(\myreg/Reg[8][3] ), .Z(\myreg/_0473_ ) );
BUF_X1 \myreg/_5980_ ( .A(\myreg/Reg[9][3] ), .Z(\myreg/_0505_ ) );
BUF_X1 \myreg/_5981_ ( .A(\myreg/Reg[10][3] ), .Z(\myreg/_0057_ ) );
BUF_X1 \myreg/_5982_ ( .A(\myreg/Reg[11][3] ), .Z(\myreg/_0089_ ) );
BUF_X1 \myreg/_5983_ ( .A(\myreg/Reg[12][3] ), .Z(\myreg/_0121_ ) );
BUF_X1 \myreg/_5984_ ( .A(\myreg/Reg[13][3] ), .Z(\myreg/_0153_ ) );
BUF_X1 \myreg/_5985_ ( .A(\myreg/Reg[14][3] ), .Z(\myreg/_0185_ ) );
BUF_X1 \myreg/_5986_ ( .A(\myreg/Reg[15][3] ), .Z(\myreg/_0217_ ) );
BUF_X1 \myreg/_5987_ ( .A(\myreg/_2373_ ), .Z(\src1_raw [3] ) );
BUF_X1 \myreg/_5988_ ( .A(\myreg/Reg[0][4] ), .Z(\myreg/_0026_ ) );
BUF_X1 \myreg/_5989_ ( .A(\myreg/Reg[1][4] ), .Z(\myreg/_0250_ ) );
BUF_X1 \myreg/_5990_ ( .A(\myreg/Reg[2][4] ), .Z(\myreg/_0282_ ) );
BUF_X1 \myreg/_5991_ ( .A(\myreg/Reg[3][4] ), .Z(\myreg/_0314_ ) );
BUF_X1 \myreg/_5992_ ( .A(\myreg/Reg[4][4] ), .Z(\myreg/_0346_ ) );
BUF_X1 \myreg/_5993_ ( .A(\myreg/Reg[5][4] ), .Z(\myreg/_0378_ ) );
BUF_X1 \myreg/_5994_ ( .A(\myreg/Reg[6][4] ), .Z(\myreg/_0410_ ) );
BUF_X1 \myreg/_5995_ ( .A(\myreg/Reg[7][4] ), .Z(\myreg/_0442_ ) );
BUF_X1 \myreg/_5996_ ( .A(\myreg/Reg[8][4] ), .Z(\myreg/_0474_ ) );
BUF_X1 \myreg/_5997_ ( .A(\myreg/Reg[9][4] ), .Z(\myreg/_0506_ ) );
BUF_X1 \myreg/_5998_ ( .A(\myreg/Reg[10][4] ), .Z(\myreg/_0058_ ) );
BUF_X1 \myreg/_5999_ ( .A(\myreg/Reg[11][4] ), .Z(\myreg/_0090_ ) );
BUF_X1 \myreg/_6000_ ( .A(\myreg/Reg[12][4] ), .Z(\myreg/_0122_ ) );
BUF_X1 \myreg/_6001_ ( .A(\myreg/Reg[13][4] ), .Z(\myreg/_0154_ ) );
BUF_X1 \myreg/_6002_ ( .A(\myreg/Reg[14][4] ), .Z(\myreg/_0186_ ) );
BUF_X1 \myreg/_6003_ ( .A(\myreg/Reg[15][4] ), .Z(\myreg/_0218_ ) );
BUF_X1 \myreg/_6004_ ( .A(\myreg/_2374_ ), .Z(\src1_raw [4] ) );
BUF_X1 \myreg/_6005_ ( .A(\myreg/Reg[0][5] ), .Z(\myreg/_0027_ ) );
BUF_X1 \myreg/_6006_ ( .A(\myreg/Reg[1][5] ), .Z(\myreg/_0251_ ) );
BUF_X1 \myreg/_6007_ ( .A(\myreg/Reg[2][5] ), .Z(\myreg/_0283_ ) );
BUF_X1 \myreg/_6008_ ( .A(\myreg/Reg[3][5] ), .Z(\myreg/_0315_ ) );
BUF_X1 \myreg/_6009_ ( .A(\myreg/Reg[4][5] ), .Z(\myreg/_0347_ ) );
BUF_X1 \myreg/_6010_ ( .A(\myreg/Reg[5][5] ), .Z(\myreg/_0379_ ) );
BUF_X1 \myreg/_6011_ ( .A(\myreg/Reg[6][5] ), .Z(\myreg/_0411_ ) );
BUF_X1 \myreg/_6012_ ( .A(\myreg/Reg[7][5] ), .Z(\myreg/_0443_ ) );
BUF_X1 \myreg/_6013_ ( .A(\myreg/Reg[8][5] ), .Z(\myreg/_0475_ ) );
BUF_X1 \myreg/_6014_ ( .A(\myreg/Reg[9][5] ), .Z(\myreg/_0507_ ) );
BUF_X1 \myreg/_6015_ ( .A(\myreg/Reg[10][5] ), .Z(\myreg/_0059_ ) );
BUF_X1 \myreg/_6016_ ( .A(\myreg/Reg[11][5] ), .Z(\myreg/_0091_ ) );
BUF_X1 \myreg/_6017_ ( .A(\myreg/Reg[12][5] ), .Z(\myreg/_0123_ ) );
BUF_X1 \myreg/_6018_ ( .A(\myreg/Reg[13][5] ), .Z(\myreg/_0155_ ) );
BUF_X1 \myreg/_6019_ ( .A(\myreg/Reg[14][5] ), .Z(\myreg/_0187_ ) );
BUF_X1 \myreg/_6020_ ( .A(\myreg/Reg[15][5] ), .Z(\myreg/_0219_ ) );
BUF_X1 \myreg/_6021_ ( .A(\myreg/_2375_ ), .Z(\src1_raw [5] ) );
BUF_X1 \myreg/_6022_ ( .A(\myreg/Reg[0][6] ), .Z(\myreg/_0028_ ) );
BUF_X1 \myreg/_6023_ ( .A(\myreg/Reg[1][6] ), .Z(\myreg/_0252_ ) );
BUF_X1 \myreg/_6024_ ( .A(\myreg/Reg[2][6] ), .Z(\myreg/_0284_ ) );
BUF_X1 \myreg/_6025_ ( .A(\myreg/Reg[3][6] ), .Z(\myreg/_0316_ ) );
BUF_X1 \myreg/_6026_ ( .A(\myreg/Reg[4][6] ), .Z(\myreg/_0348_ ) );
BUF_X1 \myreg/_6027_ ( .A(\myreg/Reg[5][6] ), .Z(\myreg/_0380_ ) );
BUF_X1 \myreg/_6028_ ( .A(\myreg/Reg[6][6] ), .Z(\myreg/_0412_ ) );
BUF_X1 \myreg/_6029_ ( .A(\myreg/Reg[7][6] ), .Z(\myreg/_0444_ ) );
BUF_X1 \myreg/_6030_ ( .A(\myreg/Reg[8][6] ), .Z(\myreg/_0476_ ) );
BUF_X1 \myreg/_6031_ ( .A(\myreg/Reg[9][6] ), .Z(\myreg/_0508_ ) );
BUF_X1 \myreg/_6032_ ( .A(\myreg/Reg[10][6] ), .Z(\myreg/_0060_ ) );
BUF_X1 \myreg/_6033_ ( .A(\myreg/Reg[11][6] ), .Z(\myreg/_0092_ ) );
BUF_X1 \myreg/_6034_ ( .A(\myreg/Reg[12][6] ), .Z(\myreg/_0124_ ) );
BUF_X1 \myreg/_6035_ ( .A(\myreg/Reg[13][6] ), .Z(\myreg/_0156_ ) );
BUF_X1 \myreg/_6036_ ( .A(\myreg/Reg[14][6] ), .Z(\myreg/_0188_ ) );
BUF_X1 \myreg/_6037_ ( .A(\myreg/Reg[15][6] ), .Z(\myreg/_0220_ ) );
BUF_X1 \myreg/_6038_ ( .A(\myreg/_2376_ ), .Z(\src1_raw [6] ) );
BUF_X1 \myreg/_6039_ ( .A(\myreg/Reg[0][7] ), .Z(\myreg/_0029_ ) );
BUF_X1 \myreg/_6040_ ( .A(\myreg/Reg[1][7] ), .Z(\myreg/_0253_ ) );
BUF_X1 \myreg/_6041_ ( .A(\myreg/Reg[2][7] ), .Z(\myreg/_0285_ ) );
BUF_X1 \myreg/_6042_ ( .A(\myreg/Reg[3][7] ), .Z(\myreg/_0317_ ) );
BUF_X1 \myreg/_6043_ ( .A(\myreg/Reg[4][7] ), .Z(\myreg/_0349_ ) );
BUF_X1 \myreg/_6044_ ( .A(\myreg/Reg[5][7] ), .Z(\myreg/_0381_ ) );
BUF_X1 \myreg/_6045_ ( .A(\myreg/Reg[6][7] ), .Z(\myreg/_0413_ ) );
BUF_X1 \myreg/_6046_ ( .A(\myreg/Reg[7][7] ), .Z(\myreg/_0445_ ) );
BUF_X1 \myreg/_6047_ ( .A(\myreg/Reg[8][7] ), .Z(\myreg/_0477_ ) );
BUF_X1 \myreg/_6048_ ( .A(\myreg/Reg[9][7] ), .Z(\myreg/_0509_ ) );
BUF_X1 \myreg/_6049_ ( .A(\myreg/Reg[10][7] ), .Z(\myreg/_0061_ ) );
BUF_X1 \myreg/_6050_ ( .A(\myreg/Reg[11][7] ), .Z(\myreg/_0093_ ) );
BUF_X1 \myreg/_6051_ ( .A(\myreg/Reg[12][7] ), .Z(\myreg/_0125_ ) );
BUF_X1 \myreg/_6052_ ( .A(\myreg/Reg[13][7] ), .Z(\myreg/_0157_ ) );
BUF_X1 \myreg/_6053_ ( .A(\myreg/Reg[14][7] ), .Z(\myreg/_0189_ ) );
BUF_X1 \myreg/_6054_ ( .A(\myreg/Reg[15][7] ), .Z(\myreg/_0221_ ) );
BUF_X1 \myreg/_6055_ ( .A(\myreg/_2377_ ), .Z(\src1_raw [7] ) );
BUF_X1 \myreg/_6056_ ( .A(\myreg/Reg[0][8] ), .Z(\myreg/_0030_ ) );
BUF_X1 \myreg/_6057_ ( .A(\myreg/Reg[1][8] ), .Z(\myreg/_0254_ ) );
BUF_X1 \myreg/_6058_ ( .A(\myreg/Reg[2][8] ), .Z(\myreg/_0286_ ) );
BUF_X1 \myreg/_6059_ ( .A(\myreg/Reg[3][8] ), .Z(\myreg/_0318_ ) );
BUF_X1 \myreg/_6060_ ( .A(\myreg/Reg[4][8] ), .Z(\myreg/_0350_ ) );
BUF_X1 \myreg/_6061_ ( .A(\myreg/Reg[5][8] ), .Z(\myreg/_0382_ ) );
BUF_X1 \myreg/_6062_ ( .A(\myreg/Reg[6][8] ), .Z(\myreg/_0414_ ) );
BUF_X1 \myreg/_6063_ ( .A(\myreg/Reg[7][8] ), .Z(\myreg/_0446_ ) );
BUF_X1 \myreg/_6064_ ( .A(\myreg/Reg[8][8] ), .Z(\myreg/_0478_ ) );
BUF_X1 \myreg/_6065_ ( .A(\myreg/Reg[9][8] ), .Z(\myreg/_0510_ ) );
BUF_X1 \myreg/_6066_ ( .A(\myreg/Reg[10][8] ), .Z(\myreg/_0062_ ) );
BUF_X1 \myreg/_6067_ ( .A(\myreg/Reg[11][8] ), .Z(\myreg/_0094_ ) );
BUF_X1 \myreg/_6068_ ( .A(\myreg/Reg[12][8] ), .Z(\myreg/_0126_ ) );
BUF_X1 \myreg/_6069_ ( .A(\myreg/Reg[13][8] ), .Z(\myreg/_0158_ ) );
BUF_X1 \myreg/_6070_ ( .A(\myreg/Reg[14][8] ), .Z(\myreg/_0190_ ) );
BUF_X1 \myreg/_6071_ ( .A(\myreg/Reg[15][8] ), .Z(\myreg/_0222_ ) );
BUF_X1 \myreg/_6072_ ( .A(\myreg/_2378_ ), .Z(\src1_raw [8] ) );
BUF_X1 \myreg/_6073_ ( .A(\myreg/Reg[0][9] ), .Z(\myreg/_0031_ ) );
BUF_X1 \myreg/_6074_ ( .A(\myreg/Reg[1][9] ), .Z(\myreg/_0255_ ) );
BUF_X1 \myreg/_6075_ ( .A(\myreg/Reg[2][9] ), .Z(\myreg/_0287_ ) );
BUF_X1 \myreg/_6076_ ( .A(\myreg/Reg[3][9] ), .Z(\myreg/_0319_ ) );
BUF_X1 \myreg/_6077_ ( .A(\myreg/Reg[4][9] ), .Z(\myreg/_0351_ ) );
BUF_X1 \myreg/_6078_ ( .A(\myreg/Reg[5][9] ), .Z(\myreg/_0383_ ) );
BUF_X1 \myreg/_6079_ ( .A(\myreg/Reg[6][9] ), .Z(\myreg/_0415_ ) );
BUF_X1 \myreg/_6080_ ( .A(\myreg/Reg[7][9] ), .Z(\myreg/_0447_ ) );
BUF_X1 \myreg/_6081_ ( .A(\myreg/Reg[8][9] ), .Z(\myreg/_0479_ ) );
BUF_X1 \myreg/_6082_ ( .A(\myreg/Reg[9][9] ), .Z(\myreg/_0511_ ) );
BUF_X1 \myreg/_6083_ ( .A(\myreg/Reg[10][9] ), .Z(\myreg/_0063_ ) );
BUF_X1 \myreg/_6084_ ( .A(\myreg/Reg[11][9] ), .Z(\myreg/_0095_ ) );
BUF_X1 \myreg/_6085_ ( .A(\myreg/Reg[12][9] ), .Z(\myreg/_0127_ ) );
BUF_X1 \myreg/_6086_ ( .A(\myreg/Reg[13][9] ), .Z(\myreg/_0159_ ) );
BUF_X1 \myreg/_6087_ ( .A(\myreg/Reg[14][9] ), .Z(\myreg/_0191_ ) );
BUF_X1 \myreg/_6088_ ( .A(\myreg/Reg[15][9] ), .Z(\myreg/_0223_ ) );
BUF_X1 \myreg/_6089_ ( .A(\myreg/_2379_ ), .Z(\src1_raw [9] ) );
BUF_X1 \myreg/_6090_ ( .A(\myreg/Reg[0][10] ), .Z(\myreg/_0001_ ) );
BUF_X1 \myreg/_6091_ ( .A(\myreg/Reg[1][10] ), .Z(\myreg/_0225_ ) );
BUF_X1 \myreg/_6092_ ( .A(\myreg/Reg[2][10] ), .Z(\myreg/_0257_ ) );
BUF_X1 \myreg/_6093_ ( .A(\myreg/Reg[3][10] ), .Z(\myreg/_0289_ ) );
BUF_X1 \myreg/_6094_ ( .A(\myreg/Reg[4][10] ), .Z(\myreg/_0321_ ) );
BUF_X1 \myreg/_6095_ ( .A(\myreg/Reg[5][10] ), .Z(\myreg/_0353_ ) );
BUF_X1 \myreg/_6096_ ( .A(\myreg/Reg[6][10] ), .Z(\myreg/_0385_ ) );
BUF_X1 \myreg/_6097_ ( .A(\myreg/Reg[7][10] ), .Z(\myreg/_0417_ ) );
BUF_X1 \myreg/_6098_ ( .A(\myreg/Reg[8][10] ), .Z(\myreg/_0449_ ) );
BUF_X1 \myreg/_6099_ ( .A(\myreg/Reg[9][10] ), .Z(\myreg/_0481_ ) );
BUF_X1 \myreg/_6100_ ( .A(\myreg/Reg[10][10] ), .Z(\myreg/_0033_ ) );
BUF_X1 \myreg/_6101_ ( .A(\myreg/Reg[11][10] ), .Z(\myreg/_0065_ ) );
BUF_X1 \myreg/_6102_ ( .A(\myreg/Reg[12][10] ), .Z(\myreg/_0097_ ) );
BUF_X1 \myreg/_6103_ ( .A(\myreg/Reg[13][10] ), .Z(\myreg/_0129_ ) );
BUF_X1 \myreg/_6104_ ( .A(\myreg/Reg[14][10] ), .Z(\myreg/_0161_ ) );
BUF_X1 \myreg/_6105_ ( .A(\myreg/Reg[15][10] ), .Z(\myreg/_0193_ ) );
BUF_X1 \myreg/_6106_ ( .A(\myreg/_2349_ ), .Z(\src1_raw [10] ) );
BUF_X1 \myreg/_6107_ ( .A(\myreg/Reg[0][11] ), .Z(\myreg/_0002_ ) );
BUF_X1 \myreg/_6108_ ( .A(\myreg/Reg[1][11] ), .Z(\myreg/_0226_ ) );
BUF_X1 \myreg/_6109_ ( .A(\myreg/Reg[2][11] ), .Z(\myreg/_0258_ ) );
BUF_X1 \myreg/_6110_ ( .A(\myreg/Reg[3][11] ), .Z(\myreg/_0290_ ) );
BUF_X1 \myreg/_6111_ ( .A(\myreg/Reg[4][11] ), .Z(\myreg/_0322_ ) );
BUF_X1 \myreg/_6112_ ( .A(\myreg/Reg[5][11] ), .Z(\myreg/_0354_ ) );
BUF_X1 \myreg/_6113_ ( .A(\myreg/Reg[6][11] ), .Z(\myreg/_0386_ ) );
BUF_X1 \myreg/_6114_ ( .A(\myreg/Reg[7][11] ), .Z(\myreg/_0418_ ) );
BUF_X1 \myreg/_6115_ ( .A(\myreg/Reg[8][11] ), .Z(\myreg/_0450_ ) );
BUF_X1 \myreg/_6116_ ( .A(\myreg/Reg[9][11] ), .Z(\myreg/_0482_ ) );
BUF_X1 \myreg/_6117_ ( .A(\myreg/Reg[10][11] ), .Z(\myreg/_0034_ ) );
BUF_X1 \myreg/_6118_ ( .A(\myreg/Reg[11][11] ), .Z(\myreg/_0066_ ) );
BUF_X1 \myreg/_6119_ ( .A(\myreg/Reg[12][11] ), .Z(\myreg/_0098_ ) );
BUF_X1 \myreg/_6120_ ( .A(\myreg/Reg[13][11] ), .Z(\myreg/_0130_ ) );
BUF_X1 \myreg/_6121_ ( .A(\myreg/Reg[14][11] ), .Z(\myreg/_0162_ ) );
BUF_X1 \myreg/_6122_ ( .A(\myreg/Reg[15][11] ), .Z(\myreg/_0194_ ) );
BUF_X1 \myreg/_6123_ ( .A(\myreg/_2350_ ), .Z(\src1_raw [11] ) );
BUF_X1 \myreg/_6124_ ( .A(\myreg/Reg[0][12] ), .Z(\myreg/_0003_ ) );
BUF_X1 \myreg/_6125_ ( .A(\myreg/Reg[1][12] ), .Z(\myreg/_0227_ ) );
BUF_X1 \myreg/_6126_ ( .A(\myreg/Reg[2][12] ), .Z(\myreg/_0259_ ) );
BUF_X1 \myreg/_6127_ ( .A(\myreg/Reg[3][12] ), .Z(\myreg/_0291_ ) );
BUF_X1 \myreg/_6128_ ( .A(\myreg/Reg[4][12] ), .Z(\myreg/_0323_ ) );
BUF_X1 \myreg/_6129_ ( .A(\myreg/Reg[5][12] ), .Z(\myreg/_0355_ ) );
BUF_X1 \myreg/_6130_ ( .A(\myreg/Reg[6][12] ), .Z(\myreg/_0387_ ) );
BUF_X1 \myreg/_6131_ ( .A(\myreg/Reg[7][12] ), .Z(\myreg/_0419_ ) );
BUF_X1 \myreg/_6132_ ( .A(\myreg/Reg[8][12] ), .Z(\myreg/_0451_ ) );
BUF_X1 \myreg/_6133_ ( .A(\myreg/Reg[9][12] ), .Z(\myreg/_0483_ ) );
BUF_X1 \myreg/_6134_ ( .A(\myreg/Reg[10][12] ), .Z(\myreg/_0035_ ) );
BUF_X1 \myreg/_6135_ ( .A(\myreg/Reg[11][12] ), .Z(\myreg/_0067_ ) );
BUF_X1 \myreg/_6136_ ( .A(\myreg/Reg[12][12] ), .Z(\myreg/_0099_ ) );
BUF_X1 \myreg/_6137_ ( .A(\myreg/Reg[13][12] ), .Z(\myreg/_0131_ ) );
BUF_X1 \myreg/_6138_ ( .A(\myreg/Reg[14][12] ), .Z(\myreg/_0163_ ) );
BUF_X1 \myreg/_6139_ ( .A(\myreg/Reg[15][12] ), .Z(\myreg/_0195_ ) );
BUF_X1 \myreg/_6140_ ( .A(\myreg/_2351_ ), .Z(\src1_raw [12] ) );
BUF_X1 \myreg/_6141_ ( .A(\myreg/Reg[0][13] ), .Z(\myreg/_0004_ ) );
BUF_X1 \myreg/_6142_ ( .A(\myreg/Reg[1][13] ), .Z(\myreg/_0228_ ) );
BUF_X1 \myreg/_6143_ ( .A(\myreg/Reg[2][13] ), .Z(\myreg/_0260_ ) );
BUF_X1 \myreg/_6144_ ( .A(\myreg/Reg[3][13] ), .Z(\myreg/_0292_ ) );
BUF_X1 \myreg/_6145_ ( .A(\myreg/Reg[4][13] ), .Z(\myreg/_0324_ ) );
BUF_X1 \myreg/_6146_ ( .A(\myreg/Reg[5][13] ), .Z(\myreg/_0356_ ) );
BUF_X1 \myreg/_6147_ ( .A(\myreg/Reg[6][13] ), .Z(\myreg/_0388_ ) );
BUF_X1 \myreg/_6148_ ( .A(\myreg/Reg[7][13] ), .Z(\myreg/_0420_ ) );
BUF_X1 \myreg/_6149_ ( .A(\myreg/Reg[8][13] ), .Z(\myreg/_0452_ ) );
BUF_X1 \myreg/_6150_ ( .A(\myreg/Reg[9][13] ), .Z(\myreg/_0484_ ) );
BUF_X1 \myreg/_6151_ ( .A(\myreg/Reg[10][13] ), .Z(\myreg/_0036_ ) );
BUF_X1 \myreg/_6152_ ( .A(\myreg/Reg[11][13] ), .Z(\myreg/_0068_ ) );
BUF_X1 \myreg/_6153_ ( .A(\myreg/Reg[12][13] ), .Z(\myreg/_0100_ ) );
BUF_X1 \myreg/_6154_ ( .A(\myreg/Reg[13][13] ), .Z(\myreg/_0132_ ) );
BUF_X1 \myreg/_6155_ ( .A(\myreg/Reg[14][13] ), .Z(\myreg/_0164_ ) );
BUF_X1 \myreg/_6156_ ( .A(\myreg/Reg[15][13] ), .Z(\myreg/_0196_ ) );
BUF_X1 \myreg/_6157_ ( .A(\myreg/_2352_ ), .Z(\src1_raw [13] ) );
BUF_X1 \myreg/_6158_ ( .A(\myreg/Reg[0][14] ), .Z(\myreg/_0005_ ) );
BUF_X1 \myreg/_6159_ ( .A(\myreg/Reg[1][14] ), .Z(\myreg/_0229_ ) );
BUF_X1 \myreg/_6160_ ( .A(\myreg/Reg[2][14] ), .Z(\myreg/_0261_ ) );
BUF_X1 \myreg/_6161_ ( .A(\myreg/Reg[3][14] ), .Z(\myreg/_0293_ ) );
BUF_X1 \myreg/_6162_ ( .A(\myreg/Reg[4][14] ), .Z(\myreg/_0325_ ) );
BUF_X1 \myreg/_6163_ ( .A(\myreg/Reg[5][14] ), .Z(\myreg/_0357_ ) );
BUF_X1 \myreg/_6164_ ( .A(\myreg/Reg[6][14] ), .Z(\myreg/_0389_ ) );
BUF_X1 \myreg/_6165_ ( .A(\myreg/Reg[7][14] ), .Z(\myreg/_0421_ ) );
BUF_X1 \myreg/_6166_ ( .A(\myreg/Reg[8][14] ), .Z(\myreg/_0453_ ) );
BUF_X1 \myreg/_6167_ ( .A(\myreg/Reg[9][14] ), .Z(\myreg/_0485_ ) );
BUF_X1 \myreg/_6168_ ( .A(\myreg/Reg[10][14] ), .Z(\myreg/_0037_ ) );
BUF_X1 \myreg/_6169_ ( .A(\myreg/Reg[11][14] ), .Z(\myreg/_0069_ ) );
BUF_X1 \myreg/_6170_ ( .A(\myreg/Reg[12][14] ), .Z(\myreg/_0101_ ) );
BUF_X1 \myreg/_6171_ ( .A(\myreg/Reg[13][14] ), .Z(\myreg/_0133_ ) );
BUF_X1 \myreg/_6172_ ( .A(\myreg/Reg[14][14] ), .Z(\myreg/_0165_ ) );
BUF_X1 \myreg/_6173_ ( .A(\myreg/Reg[15][14] ), .Z(\myreg/_0197_ ) );
BUF_X1 \myreg/_6174_ ( .A(\myreg/_2353_ ), .Z(\src1_raw [14] ) );
BUF_X1 \myreg/_6175_ ( .A(\myreg/Reg[0][15] ), .Z(\myreg/_0006_ ) );
BUF_X1 \myreg/_6176_ ( .A(\myreg/Reg[1][15] ), .Z(\myreg/_0230_ ) );
BUF_X1 \myreg/_6177_ ( .A(\myreg/Reg[2][15] ), .Z(\myreg/_0262_ ) );
BUF_X1 \myreg/_6178_ ( .A(\myreg/Reg[3][15] ), .Z(\myreg/_0294_ ) );
BUF_X1 \myreg/_6179_ ( .A(\myreg/Reg[4][15] ), .Z(\myreg/_0326_ ) );
BUF_X1 \myreg/_6180_ ( .A(\myreg/Reg[5][15] ), .Z(\myreg/_0358_ ) );
BUF_X1 \myreg/_6181_ ( .A(\myreg/Reg[6][15] ), .Z(\myreg/_0390_ ) );
BUF_X1 \myreg/_6182_ ( .A(\myreg/Reg[7][15] ), .Z(\myreg/_0422_ ) );
BUF_X1 \myreg/_6183_ ( .A(\myreg/Reg[8][15] ), .Z(\myreg/_0454_ ) );
BUF_X1 \myreg/_6184_ ( .A(\myreg/Reg[9][15] ), .Z(\myreg/_0486_ ) );
BUF_X1 \myreg/_6185_ ( .A(\myreg/Reg[10][15] ), .Z(\myreg/_0038_ ) );
BUF_X1 \myreg/_6186_ ( .A(\myreg/Reg[11][15] ), .Z(\myreg/_0070_ ) );
BUF_X1 \myreg/_6187_ ( .A(\myreg/Reg[12][15] ), .Z(\myreg/_0102_ ) );
BUF_X1 \myreg/_6188_ ( .A(\myreg/Reg[13][15] ), .Z(\myreg/_0134_ ) );
BUF_X1 \myreg/_6189_ ( .A(\myreg/Reg[14][15] ), .Z(\myreg/_0166_ ) );
BUF_X1 \myreg/_6190_ ( .A(\myreg/Reg[15][15] ), .Z(\myreg/_0198_ ) );
BUF_X1 \myreg/_6191_ ( .A(\myreg/_2354_ ), .Z(\src1_raw [15] ) );
BUF_X1 \myreg/_6192_ ( .A(\myreg/Reg[0][16] ), .Z(\myreg/_0007_ ) );
BUF_X1 \myreg/_6193_ ( .A(\myreg/Reg[1][16] ), .Z(\myreg/_0231_ ) );
BUF_X1 \myreg/_6194_ ( .A(\myreg/Reg[2][16] ), .Z(\myreg/_0263_ ) );
BUF_X1 \myreg/_6195_ ( .A(\myreg/Reg[3][16] ), .Z(\myreg/_0295_ ) );
BUF_X1 \myreg/_6196_ ( .A(\myreg/Reg[4][16] ), .Z(\myreg/_0327_ ) );
BUF_X1 \myreg/_6197_ ( .A(\myreg/Reg[5][16] ), .Z(\myreg/_0359_ ) );
BUF_X1 \myreg/_6198_ ( .A(\myreg/Reg[6][16] ), .Z(\myreg/_0391_ ) );
BUF_X1 \myreg/_6199_ ( .A(\myreg/Reg[7][16] ), .Z(\myreg/_0423_ ) );
BUF_X1 \myreg/_6200_ ( .A(\myreg/Reg[8][16] ), .Z(\myreg/_0455_ ) );
BUF_X1 \myreg/_6201_ ( .A(\myreg/Reg[9][16] ), .Z(\myreg/_0487_ ) );
BUF_X1 \myreg/_6202_ ( .A(\myreg/Reg[10][16] ), .Z(\myreg/_0039_ ) );
BUF_X1 \myreg/_6203_ ( .A(\myreg/Reg[11][16] ), .Z(\myreg/_0071_ ) );
BUF_X1 \myreg/_6204_ ( .A(\myreg/Reg[12][16] ), .Z(\myreg/_0103_ ) );
BUF_X1 \myreg/_6205_ ( .A(\myreg/Reg[13][16] ), .Z(\myreg/_0135_ ) );
BUF_X1 \myreg/_6206_ ( .A(\myreg/Reg[14][16] ), .Z(\myreg/_0167_ ) );
BUF_X1 \myreg/_6207_ ( .A(\myreg/Reg[15][16] ), .Z(\myreg/_0199_ ) );
BUF_X1 \myreg/_6208_ ( .A(\myreg/_2355_ ), .Z(\src1_raw [16] ) );
BUF_X1 \myreg/_6209_ ( .A(\myreg/Reg[0][17] ), .Z(\myreg/_0008_ ) );
BUF_X1 \myreg/_6210_ ( .A(\myreg/Reg[1][17] ), .Z(\myreg/_0232_ ) );
BUF_X1 \myreg/_6211_ ( .A(\myreg/Reg[2][17] ), .Z(\myreg/_0264_ ) );
BUF_X1 \myreg/_6212_ ( .A(\myreg/Reg[3][17] ), .Z(\myreg/_0296_ ) );
BUF_X1 \myreg/_6213_ ( .A(\myreg/Reg[4][17] ), .Z(\myreg/_0328_ ) );
BUF_X1 \myreg/_6214_ ( .A(\myreg/Reg[5][17] ), .Z(\myreg/_0360_ ) );
BUF_X1 \myreg/_6215_ ( .A(\myreg/Reg[6][17] ), .Z(\myreg/_0392_ ) );
BUF_X1 \myreg/_6216_ ( .A(\myreg/Reg[7][17] ), .Z(\myreg/_0424_ ) );
BUF_X1 \myreg/_6217_ ( .A(\myreg/Reg[8][17] ), .Z(\myreg/_0456_ ) );
BUF_X1 \myreg/_6218_ ( .A(\myreg/Reg[9][17] ), .Z(\myreg/_0488_ ) );
BUF_X1 \myreg/_6219_ ( .A(\myreg/Reg[10][17] ), .Z(\myreg/_0040_ ) );
BUF_X1 \myreg/_6220_ ( .A(\myreg/Reg[11][17] ), .Z(\myreg/_0072_ ) );
BUF_X1 \myreg/_6221_ ( .A(\myreg/Reg[12][17] ), .Z(\myreg/_0104_ ) );
BUF_X1 \myreg/_6222_ ( .A(\myreg/Reg[13][17] ), .Z(\myreg/_0136_ ) );
BUF_X1 \myreg/_6223_ ( .A(\myreg/Reg[14][17] ), .Z(\myreg/_0168_ ) );
BUF_X1 \myreg/_6224_ ( .A(\myreg/Reg[15][17] ), .Z(\myreg/_0200_ ) );
BUF_X1 \myreg/_6225_ ( .A(\myreg/_2356_ ), .Z(\src1_raw [17] ) );
BUF_X1 \myreg/_6226_ ( .A(\myreg/Reg[0][18] ), .Z(\myreg/_0009_ ) );
BUF_X1 \myreg/_6227_ ( .A(\myreg/Reg[1][18] ), .Z(\myreg/_0233_ ) );
BUF_X1 \myreg/_6228_ ( .A(\myreg/Reg[2][18] ), .Z(\myreg/_0265_ ) );
BUF_X1 \myreg/_6229_ ( .A(\myreg/Reg[3][18] ), .Z(\myreg/_0297_ ) );
BUF_X1 \myreg/_6230_ ( .A(\myreg/Reg[4][18] ), .Z(\myreg/_0329_ ) );
BUF_X1 \myreg/_6231_ ( .A(\myreg/Reg[5][18] ), .Z(\myreg/_0361_ ) );
BUF_X1 \myreg/_6232_ ( .A(\myreg/Reg[6][18] ), .Z(\myreg/_0393_ ) );
BUF_X1 \myreg/_6233_ ( .A(\myreg/Reg[7][18] ), .Z(\myreg/_0425_ ) );
BUF_X1 \myreg/_6234_ ( .A(\myreg/Reg[8][18] ), .Z(\myreg/_0457_ ) );
BUF_X1 \myreg/_6235_ ( .A(\myreg/Reg[9][18] ), .Z(\myreg/_0489_ ) );
BUF_X1 \myreg/_6236_ ( .A(\myreg/Reg[10][18] ), .Z(\myreg/_0041_ ) );
BUF_X1 \myreg/_6237_ ( .A(\myreg/Reg[11][18] ), .Z(\myreg/_0073_ ) );
BUF_X1 \myreg/_6238_ ( .A(\myreg/Reg[12][18] ), .Z(\myreg/_0105_ ) );
BUF_X1 \myreg/_6239_ ( .A(\myreg/Reg[13][18] ), .Z(\myreg/_0137_ ) );
BUF_X1 \myreg/_6240_ ( .A(\myreg/Reg[14][18] ), .Z(\myreg/_0169_ ) );
BUF_X1 \myreg/_6241_ ( .A(\myreg/Reg[15][18] ), .Z(\myreg/_0201_ ) );
BUF_X1 \myreg/_6242_ ( .A(\myreg/_2357_ ), .Z(\src1_raw [18] ) );
BUF_X1 \myreg/_6243_ ( .A(\myreg/Reg[0][19] ), .Z(\myreg/_0010_ ) );
BUF_X1 \myreg/_6244_ ( .A(\myreg/Reg[1][19] ), .Z(\myreg/_0234_ ) );
BUF_X1 \myreg/_6245_ ( .A(\myreg/Reg[2][19] ), .Z(\myreg/_0266_ ) );
BUF_X1 \myreg/_6246_ ( .A(\myreg/Reg[3][19] ), .Z(\myreg/_0298_ ) );
BUF_X1 \myreg/_6247_ ( .A(\myreg/Reg[4][19] ), .Z(\myreg/_0330_ ) );
BUF_X1 \myreg/_6248_ ( .A(\myreg/Reg[5][19] ), .Z(\myreg/_0362_ ) );
BUF_X1 \myreg/_6249_ ( .A(\myreg/Reg[6][19] ), .Z(\myreg/_0394_ ) );
BUF_X1 \myreg/_6250_ ( .A(\myreg/Reg[7][19] ), .Z(\myreg/_0426_ ) );
BUF_X1 \myreg/_6251_ ( .A(\myreg/Reg[8][19] ), .Z(\myreg/_0458_ ) );
BUF_X1 \myreg/_6252_ ( .A(\myreg/Reg[9][19] ), .Z(\myreg/_0490_ ) );
BUF_X1 \myreg/_6253_ ( .A(\myreg/Reg[10][19] ), .Z(\myreg/_0042_ ) );
BUF_X1 \myreg/_6254_ ( .A(\myreg/Reg[11][19] ), .Z(\myreg/_0074_ ) );
BUF_X1 \myreg/_6255_ ( .A(\myreg/Reg[12][19] ), .Z(\myreg/_0106_ ) );
BUF_X1 \myreg/_6256_ ( .A(\myreg/Reg[13][19] ), .Z(\myreg/_0138_ ) );
BUF_X1 \myreg/_6257_ ( .A(\myreg/Reg[14][19] ), .Z(\myreg/_0170_ ) );
BUF_X1 \myreg/_6258_ ( .A(\myreg/Reg[15][19] ), .Z(\myreg/_0202_ ) );
BUF_X1 \myreg/_6259_ ( .A(\myreg/_2358_ ), .Z(\src1_raw [19] ) );
BUF_X1 \myreg/_6260_ ( .A(\myreg/Reg[0][20] ), .Z(\myreg/_0012_ ) );
BUF_X1 \myreg/_6261_ ( .A(\myreg/Reg[1][20] ), .Z(\myreg/_0236_ ) );
BUF_X1 \myreg/_6262_ ( .A(\myreg/Reg[2][20] ), .Z(\myreg/_0268_ ) );
BUF_X1 \myreg/_6263_ ( .A(\myreg/Reg[3][20] ), .Z(\myreg/_0300_ ) );
BUF_X1 \myreg/_6264_ ( .A(\myreg/Reg[4][20] ), .Z(\myreg/_0332_ ) );
BUF_X1 \myreg/_6265_ ( .A(\myreg/Reg[5][20] ), .Z(\myreg/_0364_ ) );
BUF_X1 \myreg/_6266_ ( .A(\myreg/Reg[6][20] ), .Z(\myreg/_0396_ ) );
BUF_X1 \myreg/_6267_ ( .A(\myreg/Reg[7][20] ), .Z(\myreg/_0428_ ) );
BUF_X1 \myreg/_6268_ ( .A(\myreg/Reg[8][20] ), .Z(\myreg/_0460_ ) );
BUF_X1 \myreg/_6269_ ( .A(\myreg/Reg[9][20] ), .Z(\myreg/_0492_ ) );
BUF_X1 \myreg/_6270_ ( .A(\myreg/Reg[10][20] ), .Z(\myreg/_0044_ ) );
BUF_X1 \myreg/_6271_ ( .A(\myreg/Reg[11][20] ), .Z(\myreg/_0076_ ) );
BUF_X1 \myreg/_6272_ ( .A(\myreg/Reg[12][20] ), .Z(\myreg/_0108_ ) );
BUF_X1 \myreg/_6273_ ( .A(\myreg/Reg[13][20] ), .Z(\myreg/_0140_ ) );
BUF_X1 \myreg/_6274_ ( .A(\myreg/Reg[14][20] ), .Z(\myreg/_0172_ ) );
BUF_X1 \myreg/_6275_ ( .A(\myreg/Reg[15][20] ), .Z(\myreg/_0204_ ) );
BUF_X1 \myreg/_6276_ ( .A(\myreg/_2360_ ), .Z(\src1_raw [20] ) );
BUF_X1 \myreg/_6277_ ( .A(\myreg/Reg[0][21] ), .Z(\myreg/_0013_ ) );
BUF_X1 \myreg/_6278_ ( .A(\myreg/Reg[1][21] ), .Z(\myreg/_0237_ ) );
BUF_X1 \myreg/_6279_ ( .A(\myreg/Reg[2][21] ), .Z(\myreg/_0269_ ) );
BUF_X1 \myreg/_6280_ ( .A(\myreg/Reg[3][21] ), .Z(\myreg/_0301_ ) );
BUF_X1 \myreg/_6281_ ( .A(\myreg/Reg[4][21] ), .Z(\myreg/_0333_ ) );
BUF_X1 \myreg/_6282_ ( .A(\myreg/Reg[5][21] ), .Z(\myreg/_0365_ ) );
BUF_X1 \myreg/_6283_ ( .A(\myreg/Reg[6][21] ), .Z(\myreg/_0397_ ) );
BUF_X1 \myreg/_6284_ ( .A(\myreg/Reg[7][21] ), .Z(\myreg/_0429_ ) );
BUF_X1 \myreg/_6285_ ( .A(\myreg/Reg[8][21] ), .Z(\myreg/_0461_ ) );
BUF_X1 \myreg/_6286_ ( .A(\myreg/Reg[9][21] ), .Z(\myreg/_0493_ ) );
BUF_X1 \myreg/_6287_ ( .A(\myreg/Reg[10][21] ), .Z(\myreg/_0045_ ) );
BUF_X1 \myreg/_6288_ ( .A(\myreg/Reg[11][21] ), .Z(\myreg/_0077_ ) );
BUF_X1 \myreg/_6289_ ( .A(\myreg/Reg[12][21] ), .Z(\myreg/_0109_ ) );
BUF_X1 \myreg/_6290_ ( .A(\myreg/Reg[13][21] ), .Z(\myreg/_0141_ ) );
BUF_X1 \myreg/_6291_ ( .A(\myreg/Reg[14][21] ), .Z(\myreg/_0173_ ) );
BUF_X1 \myreg/_6292_ ( .A(\myreg/Reg[15][21] ), .Z(\myreg/_0205_ ) );
BUF_X1 \myreg/_6293_ ( .A(\myreg/_2361_ ), .Z(\src1_raw [21] ) );
BUF_X1 \myreg/_6294_ ( .A(\myreg/Reg[0][22] ), .Z(\myreg/_0014_ ) );
BUF_X1 \myreg/_6295_ ( .A(\myreg/Reg[1][22] ), .Z(\myreg/_0238_ ) );
BUF_X1 \myreg/_6296_ ( .A(\myreg/Reg[2][22] ), .Z(\myreg/_0270_ ) );
BUF_X1 \myreg/_6297_ ( .A(\myreg/Reg[3][22] ), .Z(\myreg/_0302_ ) );
BUF_X1 \myreg/_6298_ ( .A(\myreg/Reg[4][22] ), .Z(\myreg/_0334_ ) );
BUF_X1 \myreg/_6299_ ( .A(\myreg/Reg[5][22] ), .Z(\myreg/_0366_ ) );
BUF_X1 \myreg/_6300_ ( .A(\myreg/Reg[6][22] ), .Z(\myreg/_0398_ ) );
BUF_X1 \myreg/_6301_ ( .A(\myreg/Reg[7][22] ), .Z(\myreg/_0430_ ) );
BUF_X1 \myreg/_6302_ ( .A(\myreg/Reg[8][22] ), .Z(\myreg/_0462_ ) );
BUF_X1 \myreg/_6303_ ( .A(\myreg/Reg[9][22] ), .Z(\myreg/_0494_ ) );
BUF_X1 \myreg/_6304_ ( .A(\myreg/Reg[10][22] ), .Z(\myreg/_0046_ ) );
BUF_X1 \myreg/_6305_ ( .A(\myreg/Reg[11][22] ), .Z(\myreg/_0078_ ) );
BUF_X1 \myreg/_6306_ ( .A(\myreg/Reg[12][22] ), .Z(\myreg/_0110_ ) );
BUF_X1 \myreg/_6307_ ( .A(\myreg/Reg[13][22] ), .Z(\myreg/_0142_ ) );
BUF_X1 \myreg/_6308_ ( .A(\myreg/Reg[14][22] ), .Z(\myreg/_0174_ ) );
BUF_X1 \myreg/_6309_ ( .A(\myreg/Reg[15][22] ), .Z(\myreg/_0206_ ) );
BUF_X1 \myreg/_6310_ ( .A(\myreg/_2362_ ), .Z(\src1_raw [22] ) );
BUF_X1 \myreg/_6311_ ( .A(\myreg/Reg[0][23] ), .Z(\myreg/_0015_ ) );
BUF_X1 \myreg/_6312_ ( .A(\myreg/Reg[1][23] ), .Z(\myreg/_0239_ ) );
BUF_X1 \myreg/_6313_ ( .A(\myreg/Reg[2][23] ), .Z(\myreg/_0271_ ) );
BUF_X1 \myreg/_6314_ ( .A(\myreg/Reg[3][23] ), .Z(\myreg/_0303_ ) );
BUF_X1 \myreg/_6315_ ( .A(\myreg/Reg[4][23] ), .Z(\myreg/_0335_ ) );
BUF_X1 \myreg/_6316_ ( .A(\myreg/Reg[5][23] ), .Z(\myreg/_0367_ ) );
BUF_X1 \myreg/_6317_ ( .A(\myreg/Reg[6][23] ), .Z(\myreg/_0399_ ) );
BUF_X1 \myreg/_6318_ ( .A(\myreg/Reg[7][23] ), .Z(\myreg/_0431_ ) );
BUF_X1 \myreg/_6319_ ( .A(\myreg/Reg[8][23] ), .Z(\myreg/_0463_ ) );
BUF_X1 \myreg/_6320_ ( .A(\myreg/Reg[9][23] ), .Z(\myreg/_0495_ ) );
BUF_X1 \myreg/_6321_ ( .A(\myreg/Reg[10][23] ), .Z(\myreg/_0047_ ) );
BUF_X1 \myreg/_6322_ ( .A(\myreg/Reg[11][23] ), .Z(\myreg/_0079_ ) );
BUF_X1 \myreg/_6323_ ( .A(\myreg/Reg[12][23] ), .Z(\myreg/_0111_ ) );
BUF_X1 \myreg/_6324_ ( .A(\myreg/Reg[13][23] ), .Z(\myreg/_0143_ ) );
BUF_X1 \myreg/_6325_ ( .A(\myreg/Reg[14][23] ), .Z(\myreg/_0175_ ) );
BUF_X1 \myreg/_6326_ ( .A(\myreg/Reg[15][23] ), .Z(\myreg/_0207_ ) );
BUF_X1 \myreg/_6327_ ( .A(\myreg/_2363_ ), .Z(\src1_raw [23] ) );
BUF_X1 \myreg/_6328_ ( .A(\myreg/Reg[0][24] ), .Z(\myreg/_0016_ ) );
BUF_X1 \myreg/_6329_ ( .A(\myreg/Reg[1][24] ), .Z(\myreg/_0240_ ) );
BUF_X1 \myreg/_6330_ ( .A(\myreg/Reg[2][24] ), .Z(\myreg/_0272_ ) );
BUF_X1 \myreg/_6331_ ( .A(\myreg/Reg[3][24] ), .Z(\myreg/_0304_ ) );
BUF_X1 \myreg/_6332_ ( .A(\myreg/Reg[4][24] ), .Z(\myreg/_0336_ ) );
BUF_X1 \myreg/_6333_ ( .A(\myreg/Reg[5][24] ), .Z(\myreg/_0368_ ) );
BUF_X1 \myreg/_6334_ ( .A(\myreg/Reg[6][24] ), .Z(\myreg/_0400_ ) );
BUF_X1 \myreg/_6335_ ( .A(\myreg/Reg[7][24] ), .Z(\myreg/_0432_ ) );
BUF_X1 \myreg/_6336_ ( .A(\myreg/Reg[8][24] ), .Z(\myreg/_0464_ ) );
BUF_X1 \myreg/_6337_ ( .A(\myreg/Reg[9][24] ), .Z(\myreg/_0496_ ) );
BUF_X1 \myreg/_6338_ ( .A(\myreg/Reg[10][24] ), .Z(\myreg/_0048_ ) );
BUF_X1 \myreg/_6339_ ( .A(\myreg/Reg[11][24] ), .Z(\myreg/_0080_ ) );
BUF_X1 \myreg/_6340_ ( .A(\myreg/Reg[12][24] ), .Z(\myreg/_0112_ ) );
BUF_X1 \myreg/_6341_ ( .A(\myreg/Reg[13][24] ), .Z(\myreg/_0144_ ) );
BUF_X1 \myreg/_6342_ ( .A(\myreg/Reg[14][24] ), .Z(\myreg/_0176_ ) );
BUF_X1 \myreg/_6343_ ( .A(\myreg/Reg[15][24] ), .Z(\myreg/_0208_ ) );
BUF_X1 \myreg/_6344_ ( .A(\myreg/_2364_ ), .Z(\src1_raw [24] ) );
BUF_X1 \myreg/_6345_ ( .A(\myreg/Reg[0][25] ), .Z(\myreg/_0017_ ) );
BUF_X1 \myreg/_6346_ ( .A(\myreg/Reg[1][25] ), .Z(\myreg/_0241_ ) );
BUF_X1 \myreg/_6347_ ( .A(\myreg/Reg[2][25] ), .Z(\myreg/_0273_ ) );
BUF_X1 \myreg/_6348_ ( .A(\myreg/Reg[3][25] ), .Z(\myreg/_0305_ ) );
BUF_X1 \myreg/_6349_ ( .A(\myreg/Reg[4][25] ), .Z(\myreg/_0337_ ) );
BUF_X1 \myreg/_6350_ ( .A(\myreg/Reg[5][25] ), .Z(\myreg/_0369_ ) );
BUF_X1 \myreg/_6351_ ( .A(\myreg/Reg[6][25] ), .Z(\myreg/_0401_ ) );
BUF_X1 \myreg/_6352_ ( .A(\myreg/Reg[7][25] ), .Z(\myreg/_0433_ ) );
BUF_X1 \myreg/_6353_ ( .A(\myreg/Reg[8][25] ), .Z(\myreg/_0465_ ) );
BUF_X1 \myreg/_6354_ ( .A(\myreg/Reg[9][25] ), .Z(\myreg/_0497_ ) );
BUF_X1 \myreg/_6355_ ( .A(\myreg/Reg[10][25] ), .Z(\myreg/_0049_ ) );
BUF_X1 \myreg/_6356_ ( .A(\myreg/Reg[11][25] ), .Z(\myreg/_0081_ ) );
BUF_X1 \myreg/_6357_ ( .A(\myreg/Reg[12][25] ), .Z(\myreg/_0113_ ) );
BUF_X1 \myreg/_6358_ ( .A(\myreg/Reg[13][25] ), .Z(\myreg/_0145_ ) );
BUF_X1 \myreg/_6359_ ( .A(\myreg/Reg[14][25] ), .Z(\myreg/_0177_ ) );
BUF_X1 \myreg/_6360_ ( .A(\myreg/Reg[15][25] ), .Z(\myreg/_0209_ ) );
BUF_X1 \myreg/_6361_ ( .A(\myreg/_2365_ ), .Z(\src1_raw [25] ) );
BUF_X1 \myreg/_6362_ ( .A(\myreg/Reg[0][26] ), .Z(\myreg/_0018_ ) );
BUF_X1 \myreg/_6363_ ( .A(\myreg/Reg[1][26] ), .Z(\myreg/_0242_ ) );
BUF_X1 \myreg/_6364_ ( .A(\myreg/Reg[2][26] ), .Z(\myreg/_0274_ ) );
BUF_X1 \myreg/_6365_ ( .A(\myreg/Reg[3][26] ), .Z(\myreg/_0306_ ) );
BUF_X1 \myreg/_6366_ ( .A(\myreg/Reg[4][26] ), .Z(\myreg/_0338_ ) );
BUF_X1 \myreg/_6367_ ( .A(\myreg/Reg[5][26] ), .Z(\myreg/_0370_ ) );
BUF_X1 \myreg/_6368_ ( .A(\myreg/Reg[6][26] ), .Z(\myreg/_0402_ ) );
BUF_X1 \myreg/_6369_ ( .A(\myreg/Reg[7][26] ), .Z(\myreg/_0434_ ) );
BUF_X1 \myreg/_6370_ ( .A(\myreg/Reg[8][26] ), .Z(\myreg/_0466_ ) );
BUF_X1 \myreg/_6371_ ( .A(\myreg/Reg[9][26] ), .Z(\myreg/_0498_ ) );
BUF_X1 \myreg/_6372_ ( .A(\myreg/Reg[10][26] ), .Z(\myreg/_0050_ ) );
BUF_X1 \myreg/_6373_ ( .A(\myreg/Reg[11][26] ), .Z(\myreg/_0082_ ) );
BUF_X1 \myreg/_6374_ ( .A(\myreg/Reg[12][26] ), .Z(\myreg/_0114_ ) );
BUF_X1 \myreg/_6375_ ( .A(\myreg/Reg[13][26] ), .Z(\myreg/_0146_ ) );
BUF_X1 \myreg/_6376_ ( .A(\myreg/Reg[14][26] ), .Z(\myreg/_0178_ ) );
BUF_X1 \myreg/_6377_ ( .A(\myreg/Reg[15][26] ), .Z(\myreg/_0210_ ) );
BUF_X1 \myreg/_6378_ ( .A(\myreg/_2366_ ), .Z(\src1_raw [26] ) );
BUF_X1 \myreg/_6379_ ( .A(\myreg/Reg[0][27] ), .Z(\myreg/_0019_ ) );
BUF_X1 \myreg/_6380_ ( .A(\myreg/Reg[1][27] ), .Z(\myreg/_0243_ ) );
BUF_X1 \myreg/_6381_ ( .A(\myreg/Reg[2][27] ), .Z(\myreg/_0275_ ) );
BUF_X1 \myreg/_6382_ ( .A(\myreg/Reg[3][27] ), .Z(\myreg/_0307_ ) );
BUF_X1 \myreg/_6383_ ( .A(\myreg/Reg[4][27] ), .Z(\myreg/_0339_ ) );
BUF_X1 \myreg/_6384_ ( .A(\myreg/Reg[5][27] ), .Z(\myreg/_0371_ ) );
BUF_X1 \myreg/_6385_ ( .A(\myreg/Reg[6][27] ), .Z(\myreg/_0403_ ) );
BUF_X1 \myreg/_6386_ ( .A(\myreg/Reg[7][27] ), .Z(\myreg/_0435_ ) );
BUF_X1 \myreg/_6387_ ( .A(\myreg/Reg[8][27] ), .Z(\myreg/_0467_ ) );
BUF_X1 \myreg/_6388_ ( .A(\myreg/Reg[9][27] ), .Z(\myreg/_0499_ ) );
BUF_X1 \myreg/_6389_ ( .A(\myreg/Reg[10][27] ), .Z(\myreg/_0051_ ) );
BUF_X1 \myreg/_6390_ ( .A(\myreg/Reg[11][27] ), .Z(\myreg/_0083_ ) );
BUF_X1 \myreg/_6391_ ( .A(\myreg/Reg[12][27] ), .Z(\myreg/_0115_ ) );
BUF_X1 \myreg/_6392_ ( .A(\myreg/Reg[13][27] ), .Z(\myreg/_0147_ ) );
BUF_X1 \myreg/_6393_ ( .A(\myreg/Reg[14][27] ), .Z(\myreg/_0179_ ) );
BUF_X1 \myreg/_6394_ ( .A(\myreg/Reg[15][27] ), .Z(\myreg/_0211_ ) );
BUF_X1 \myreg/_6395_ ( .A(\myreg/_2367_ ), .Z(\src1_raw [27] ) );
BUF_X1 \myreg/_6396_ ( .A(\myreg/Reg[0][28] ), .Z(\myreg/_0020_ ) );
BUF_X1 \myreg/_6397_ ( .A(\myreg/Reg[1][28] ), .Z(\myreg/_0244_ ) );
BUF_X1 \myreg/_6398_ ( .A(\myreg/Reg[2][28] ), .Z(\myreg/_0276_ ) );
BUF_X1 \myreg/_6399_ ( .A(\myreg/Reg[3][28] ), .Z(\myreg/_0308_ ) );
BUF_X1 \myreg/_6400_ ( .A(\myreg/Reg[4][28] ), .Z(\myreg/_0340_ ) );
BUF_X1 \myreg/_6401_ ( .A(\myreg/Reg[5][28] ), .Z(\myreg/_0372_ ) );
BUF_X1 \myreg/_6402_ ( .A(\myreg/Reg[6][28] ), .Z(\myreg/_0404_ ) );
BUF_X1 \myreg/_6403_ ( .A(\myreg/Reg[7][28] ), .Z(\myreg/_0436_ ) );
BUF_X1 \myreg/_6404_ ( .A(\myreg/Reg[8][28] ), .Z(\myreg/_0468_ ) );
BUF_X1 \myreg/_6405_ ( .A(\myreg/Reg[9][28] ), .Z(\myreg/_0500_ ) );
BUF_X1 \myreg/_6406_ ( .A(\myreg/Reg[10][28] ), .Z(\myreg/_0052_ ) );
BUF_X1 \myreg/_6407_ ( .A(\myreg/Reg[11][28] ), .Z(\myreg/_0084_ ) );
BUF_X1 \myreg/_6408_ ( .A(\myreg/Reg[12][28] ), .Z(\myreg/_0116_ ) );
BUF_X1 \myreg/_6409_ ( .A(\myreg/Reg[13][28] ), .Z(\myreg/_0148_ ) );
BUF_X1 \myreg/_6410_ ( .A(\myreg/Reg[14][28] ), .Z(\myreg/_0180_ ) );
BUF_X1 \myreg/_6411_ ( .A(\myreg/Reg[15][28] ), .Z(\myreg/_0212_ ) );
BUF_X1 \myreg/_6412_ ( .A(\myreg/_2368_ ), .Z(\src1_raw [28] ) );
BUF_X1 \myreg/_6413_ ( .A(\myreg/Reg[0][29] ), .Z(\myreg/_0021_ ) );
BUF_X1 \myreg/_6414_ ( .A(\myreg/Reg[1][29] ), .Z(\myreg/_0245_ ) );
BUF_X1 \myreg/_6415_ ( .A(\myreg/Reg[2][29] ), .Z(\myreg/_0277_ ) );
BUF_X1 \myreg/_6416_ ( .A(\myreg/Reg[3][29] ), .Z(\myreg/_0309_ ) );
BUF_X1 \myreg/_6417_ ( .A(\myreg/Reg[4][29] ), .Z(\myreg/_0341_ ) );
BUF_X1 \myreg/_6418_ ( .A(\myreg/Reg[5][29] ), .Z(\myreg/_0373_ ) );
BUF_X1 \myreg/_6419_ ( .A(\myreg/Reg[6][29] ), .Z(\myreg/_0405_ ) );
BUF_X1 \myreg/_6420_ ( .A(\myreg/Reg[7][29] ), .Z(\myreg/_0437_ ) );
BUF_X1 \myreg/_6421_ ( .A(\myreg/Reg[8][29] ), .Z(\myreg/_0469_ ) );
BUF_X1 \myreg/_6422_ ( .A(\myreg/Reg[9][29] ), .Z(\myreg/_0501_ ) );
BUF_X1 \myreg/_6423_ ( .A(\myreg/Reg[10][29] ), .Z(\myreg/_0053_ ) );
BUF_X1 \myreg/_6424_ ( .A(\myreg/Reg[11][29] ), .Z(\myreg/_0085_ ) );
BUF_X1 \myreg/_6425_ ( .A(\myreg/Reg[12][29] ), .Z(\myreg/_0117_ ) );
BUF_X1 \myreg/_6426_ ( .A(\myreg/Reg[13][29] ), .Z(\myreg/_0149_ ) );
BUF_X1 \myreg/_6427_ ( .A(\myreg/Reg[14][29] ), .Z(\myreg/_0181_ ) );
BUF_X1 \myreg/_6428_ ( .A(\myreg/Reg[15][29] ), .Z(\myreg/_0213_ ) );
BUF_X1 \myreg/_6429_ ( .A(\myreg/_2369_ ), .Z(\src1_raw [29] ) );
BUF_X1 \myreg/_6430_ ( .A(\myreg/Reg[0][30] ), .Z(\myreg/_0023_ ) );
BUF_X1 \myreg/_6431_ ( .A(\myreg/Reg[1][30] ), .Z(\myreg/_0247_ ) );
BUF_X1 \myreg/_6432_ ( .A(\myreg/Reg[2][30] ), .Z(\myreg/_0279_ ) );
BUF_X1 \myreg/_6433_ ( .A(\myreg/Reg[3][30] ), .Z(\myreg/_0311_ ) );
BUF_X1 \myreg/_6434_ ( .A(\myreg/Reg[4][30] ), .Z(\myreg/_0343_ ) );
BUF_X1 \myreg/_6435_ ( .A(\myreg/Reg[5][30] ), .Z(\myreg/_0375_ ) );
BUF_X1 \myreg/_6436_ ( .A(\myreg/Reg[6][30] ), .Z(\myreg/_0407_ ) );
BUF_X1 \myreg/_6437_ ( .A(\myreg/Reg[7][30] ), .Z(\myreg/_0439_ ) );
BUF_X1 \myreg/_6438_ ( .A(\myreg/Reg[8][30] ), .Z(\myreg/_0471_ ) );
BUF_X1 \myreg/_6439_ ( .A(\myreg/Reg[9][30] ), .Z(\myreg/_0503_ ) );
BUF_X1 \myreg/_6440_ ( .A(\myreg/Reg[10][30] ), .Z(\myreg/_0055_ ) );
BUF_X1 \myreg/_6441_ ( .A(\myreg/Reg[11][30] ), .Z(\myreg/_0087_ ) );
BUF_X1 \myreg/_6442_ ( .A(\myreg/Reg[12][30] ), .Z(\myreg/_0119_ ) );
BUF_X1 \myreg/_6443_ ( .A(\myreg/Reg[13][30] ), .Z(\myreg/_0151_ ) );
BUF_X1 \myreg/_6444_ ( .A(\myreg/Reg[14][30] ), .Z(\myreg/_0183_ ) );
BUF_X1 \myreg/_6445_ ( .A(\myreg/Reg[15][30] ), .Z(\myreg/_0215_ ) );
BUF_X1 \myreg/_6446_ ( .A(\myreg/_2371_ ), .Z(\src1_raw [30] ) );
BUF_X1 \myreg/_6447_ ( .A(\myreg/Reg[0][31] ), .Z(\myreg/_0024_ ) );
BUF_X1 \myreg/_6448_ ( .A(\myreg/Reg[1][31] ), .Z(\myreg/_0248_ ) );
BUF_X1 \myreg/_6449_ ( .A(\myreg/Reg[2][31] ), .Z(\myreg/_0280_ ) );
BUF_X1 \myreg/_6450_ ( .A(\myreg/Reg[3][31] ), .Z(\myreg/_0312_ ) );
BUF_X1 \myreg/_6451_ ( .A(\myreg/Reg[4][31] ), .Z(\myreg/_0344_ ) );
BUF_X1 \myreg/_6452_ ( .A(\myreg/Reg[5][31] ), .Z(\myreg/_0376_ ) );
BUF_X1 \myreg/_6453_ ( .A(\myreg/Reg[6][31] ), .Z(\myreg/_0408_ ) );
BUF_X1 \myreg/_6454_ ( .A(\myreg/Reg[7][31] ), .Z(\myreg/_0440_ ) );
BUF_X1 \myreg/_6455_ ( .A(\myreg/Reg[8][31] ), .Z(\myreg/_0472_ ) );
BUF_X1 \myreg/_6456_ ( .A(\myreg/Reg[9][31] ), .Z(\myreg/_0504_ ) );
BUF_X1 \myreg/_6457_ ( .A(\myreg/Reg[10][31] ), .Z(\myreg/_0056_ ) );
BUF_X1 \myreg/_6458_ ( .A(\myreg/Reg[11][31] ), .Z(\myreg/_0088_ ) );
BUF_X1 \myreg/_6459_ ( .A(\myreg/Reg[12][31] ), .Z(\myreg/_0120_ ) );
BUF_X1 \myreg/_6460_ ( .A(\myreg/Reg[13][31] ), .Z(\myreg/_0152_ ) );
BUF_X1 \myreg/_6461_ ( .A(\myreg/Reg[14][31] ), .Z(\myreg/_0184_ ) );
BUF_X1 \myreg/_6462_ ( .A(\myreg/Reg[15][31] ), .Z(\myreg/_0216_ ) );
BUF_X1 \myreg/_6463_ ( .A(\myreg/_2372_ ), .Z(\src1_raw [31] ) );
BUF_X1 \myreg/_6464_ ( .A(\ID_EX_rs2 [0] ), .Z(\myreg/_2344_ ) );
BUF_X1 \myreg/_6465_ ( .A(\ID_EX_rs2 [1] ), .Z(\myreg/_2345_ ) );
BUF_X1 \myreg/_6466_ ( .A(\ID_EX_rs2 [2] ), .Z(\myreg/_2346_ ) );
BUF_X1 \myreg/_6467_ ( .A(\ID_EX_rs2 [3] ), .Z(\myreg/_2347_ ) );
BUF_X1 \myreg/_6468_ ( .A(\myreg/_2380_ ), .Z(\src2_raw [0] ) );
BUF_X1 \myreg/_6469_ ( .A(\myreg/_2391_ ), .Z(\src2_raw [1] ) );
BUF_X1 \myreg/_6470_ ( .A(\myreg/_2402_ ), .Z(\src2_raw [2] ) );
BUF_X1 \myreg/_6471_ ( .A(\myreg/_2405_ ), .Z(\src2_raw [3] ) );
BUF_X1 \myreg/_6472_ ( .A(\myreg/_2406_ ), .Z(\src2_raw [4] ) );
BUF_X1 \myreg/_6473_ ( .A(\myreg/_2407_ ), .Z(\src2_raw [5] ) );
BUF_X1 \myreg/_6474_ ( .A(\myreg/_2408_ ), .Z(\src2_raw [6] ) );
BUF_X1 \myreg/_6475_ ( .A(\myreg/_2409_ ), .Z(\src2_raw [7] ) );
BUF_X1 \myreg/_6476_ ( .A(\myreg/_2410_ ), .Z(\src2_raw [8] ) );
BUF_X1 \myreg/_6477_ ( .A(\myreg/_2411_ ), .Z(\src2_raw [9] ) );
BUF_X1 \myreg/_6478_ ( .A(\myreg/_2381_ ), .Z(\src2_raw [10] ) );
BUF_X1 \myreg/_6479_ ( .A(\myreg/_2382_ ), .Z(\src2_raw [11] ) );
BUF_X1 \myreg/_6480_ ( .A(\myreg/_2383_ ), .Z(\src2_raw [12] ) );
BUF_X1 \myreg/_6481_ ( .A(\myreg/_2384_ ), .Z(\src2_raw [13] ) );
BUF_X1 \myreg/_6482_ ( .A(\myreg/_2385_ ), .Z(\src2_raw [14] ) );
BUF_X1 \myreg/_6483_ ( .A(\myreg/_2386_ ), .Z(\src2_raw [15] ) );
BUF_X1 \myreg/_6484_ ( .A(\myreg/_2387_ ), .Z(\src2_raw [16] ) );
BUF_X1 \myreg/_6485_ ( .A(\myreg/_2388_ ), .Z(\src2_raw [17] ) );
BUF_X1 \myreg/_6486_ ( .A(\myreg/_2389_ ), .Z(\src2_raw [18] ) );
BUF_X1 \myreg/_6487_ ( .A(\myreg/_2390_ ), .Z(\src2_raw [19] ) );
BUF_X1 \myreg/_6488_ ( .A(\myreg/_2392_ ), .Z(\src2_raw [20] ) );
BUF_X1 \myreg/_6489_ ( .A(\myreg/_2393_ ), .Z(\src2_raw [21] ) );
BUF_X1 \myreg/_6490_ ( .A(\myreg/_2394_ ), .Z(\src2_raw [22] ) );
BUF_X1 \myreg/_6491_ ( .A(\myreg/_2395_ ), .Z(\src2_raw [23] ) );
BUF_X1 \myreg/_6492_ ( .A(\myreg/_2396_ ), .Z(\src2_raw [24] ) );
BUF_X1 \myreg/_6493_ ( .A(\myreg/_2397_ ), .Z(\src2_raw [25] ) );
BUF_X1 \myreg/_6494_ ( .A(\myreg/_2398_ ), .Z(\src2_raw [26] ) );
BUF_X1 \myreg/_6495_ ( .A(\myreg/_2399_ ), .Z(\src2_raw [27] ) );
BUF_X1 \myreg/_6496_ ( .A(\myreg/_2400_ ), .Z(\src2_raw [28] ) );
BUF_X1 \myreg/_6497_ ( .A(\myreg/_2401_ ), .Z(\src2_raw [29] ) );
BUF_X1 \myreg/_6498_ ( .A(\myreg/_2403_ ), .Z(\src2_raw [30] ) );
BUF_X1 \myreg/_6499_ ( .A(\myreg/_2404_ ), .Z(\src2_raw [31] ) );
BUF_X1 \myreg/_6500_ ( .A(\myreg/_0512_ ), .Z(\myreg/_2962_ ) );
BUF_X1 \myreg/_6501_ ( .A(\myreg/_0513_ ), .Z(\myreg/_2963_ ) );
BUF_X1 \myreg/_6502_ ( .A(\myreg/_0514_ ), .Z(\myreg/_2964_ ) );
BUF_X1 \myreg/_6503_ ( .A(\myreg/_0515_ ), .Z(\myreg/_2965_ ) );
BUF_X1 \myreg/_6504_ ( .A(\myreg/_0516_ ), .Z(\myreg/_2966_ ) );
BUF_X1 \myreg/_6505_ ( .A(\myreg/_0517_ ), .Z(\myreg/_2967_ ) );
BUF_X1 \myreg/_6506_ ( .A(\myreg/_0518_ ), .Z(\myreg/_2968_ ) );
BUF_X1 \myreg/_6507_ ( .A(\myreg/_0519_ ), .Z(\myreg/_2969_ ) );
BUF_X1 \myreg/_6508_ ( .A(\myreg/_0520_ ), .Z(\myreg/_2970_ ) );
BUF_X1 \myreg/_6509_ ( .A(\myreg/_0521_ ), .Z(\myreg/_2971_ ) );
BUF_X1 \myreg/_6510_ ( .A(\myreg/_0522_ ), .Z(\myreg/_2972_ ) );
BUF_X1 \myreg/_6511_ ( .A(\myreg/_0523_ ), .Z(\myreg/_2973_ ) );
BUF_X1 \myreg/_6512_ ( .A(\myreg/_0524_ ), .Z(\myreg/_2974_ ) );
BUF_X1 \myreg/_6513_ ( .A(\myreg/_0525_ ), .Z(\myreg/_2975_ ) );
BUF_X1 \myreg/_6514_ ( .A(\myreg/_0526_ ), .Z(\myreg/_2976_ ) );
BUF_X1 \myreg/_6515_ ( .A(\myreg/_0527_ ), .Z(\myreg/_2977_ ) );
BUF_X1 \myreg/_6516_ ( .A(\myreg/_0528_ ), .Z(\myreg/_2978_ ) );
BUF_X1 \myreg/_6517_ ( .A(\myreg/_0529_ ), .Z(\myreg/_2979_ ) );
BUF_X1 \myreg/_6518_ ( .A(\myreg/_0530_ ), .Z(\myreg/_2980_ ) );
BUF_X1 \myreg/_6519_ ( .A(\myreg/_0531_ ), .Z(\myreg/_2981_ ) );
BUF_X1 \myreg/_6520_ ( .A(\myreg/_0532_ ), .Z(\myreg/_2982_ ) );
BUF_X1 \myreg/_6521_ ( .A(\myreg/_0533_ ), .Z(\myreg/_2983_ ) );
BUF_X1 \myreg/_6522_ ( .A(\myreg/_0534_ ), .Z(\myreg/_2984_ ) );
BUF_X1 \myreg/_6523_ ( .A(\myreg/_0535_ ), .Z(\myreg/_2985_ ) );
BUF_X1 \myreg/_6524_ ( .A(\myreg/_0536_ ), .Z(\myreg/_2986_ ) );
BUF_X1 \myreg/_6525_ ( .A(\myreg/_0537_ ), .Z(\myreg/_2987_ ) );
BUF_X1 \myreg/_6526_ ( .A(\myreg/_0538_ ), .Z(\myreg/_2988_ ) );
BUF_X1 \myreg/_6527_ ( .A(\myreg/_0539_ ), .Z(\myreg/_2989_ ) );
BUF_X1 \myreg/_6528_ ( .A(\myreg/_0540_ ), .Z(\myreg/_2990_ ) );
BUF_X1 \myreg/_6529_ ( .A(\myreg/_0541_ ), .Z(\myreg/_2991_ ) );
BUF_X1 \myreg/_6530_ ( .A(\myreg/_0542_ ), .Z(\myreg/_2992_ ) );
BUF_X1 \myreg/_6531_ ( .A(\myreg/_0543_ ), .Z(\myreg/_2993_ ) );
BUF_X1 \myreg/_6532_ ( .A(\myreg/_0544_ ), .Z(\myreg/_2994_ ) );
BUF_X1 \myreg/_6533_ ( .A(\myreg/_0545_ ), .Z(\myreg/_2995_ ) );
BUF_X1 \myreg/_6534_ ( .A(\myreg/_0546_ ), .Z(\myreg/_2996_ ) );
BUF_X1 \myreg/_6535_ ( .A(\myreg/_0547_ ), .Z(\myreg/_2997_ ) );
BUF_X1 \myreg/_6536_ ( .A(\myreg/_0548_ ), .Z(\myreg/_2998_ ) );
BUF_X1 \myreg/_6537_ ( .A(\myreg/_0549_ ), .Z(\myreg/_2999_ ) );
BUF_X1 \myreg/_6538_ ( .A(\myreg/_0550_ ), .Z(\myreg/_3000_ ) );
BUF_X1 \myreg/_6539_ ( .A(\myreg/_0551_ ), .Z(\myreg/_3001_ ) );
BUF_X1 \myreg/_6540_ ( .A(\myreg/_0552_ ), .Z(\myreg/_3002_ ) );
BUF_X1 \myreg/_6541_ ( .A(\myreg/_0553_ ), .Z(\myreg/_3003_ ) );
BUF_X1 \myreg/_6542_ ( .A(\myreg/_0554_ ), .Z(\myreg/_3004_ ) );
BUF_X1 \myreg/_6543_ ( .A(\myreg/_0555_ ), .Z(\myreg/_3005_ ) );
BUF_X1 \myreg/_6544_ ( .A(\myreg/_0556_ ), .Z(\myreg/_3006_ ) );
BUF_X1 \myreg/_6545_ ( .A(\myreg/_0557_ ), .Z(\myreg/_3007_ ) );
BUF_X1 \myreg/_6546_ ( .A(\myreg/_0558_ ), .Z(\myreg/_3008_ ) );
BUF_X1 \myreg/_6547_ ( .A(\myreg/_0559_ ), .Z(\myreg/_3009_ ) );
BUF_X1 \myreg/_6548_ ( .A(\myreg/_0560_ ), .Z(\myreg/_3010_ ) );
BUF_X1 \myreg/_6549_ ( .A(\myreg/_0561_ ), .Z(\myreg/_3011_ ) );
BUF_X1 \myreg/_6550_ ( .A(\myreg/_0562_ ), .Z(\myreg/_3012_ ) );
BUF_X1 \myreg/_6551_ ( .A(\myreg/_0563_ ), .Z(\myreg/_3013_ ) );
BUF_X1 \myreg/_6552_ ( .A(\myreg/_0564_ ), .Z(\myreg/_3014_ ) );
BUF_X1 \myreg/_6553_ ( .A(\myreg/_0565_ ), .Z(\myreg/_3015_ ) );
BUF_X1 \myreg/_6554_ ( .A(\myreg/_0566_ ), .Z(\myreg/_3016_ ) );
BUF_X1 \myreg/_6555_ ( .A(\myreg/_0567_ ), .Z(\myreg/_3017_ ) );
BUF_X1 \myreg/_6556_ ( .A(\myreg/_0568_ ), .Z(\myreg/_3018_ ) );
BUF_X1 \myreg/_6557_ ( .A(\myreg/_0569_ ), .Z(\myreg/_3019_ ) );
BUF_X1 \myreg/_6558_ ( .A(\myreg/_0570_ ), .Z(\myreg/_3020_ ) );
BUF_X1 \myreg/_6559_ ( .A(\myreg/_0571_ ), .Z(\myreg/_3021_ ) );
BUF_X1 \myreg/_6560_ ( .A(\myreg/_0572_ ), .Z(\myreg/_3022_ ) );
BUF_X1 \myreg/_6561_ ( .A(\myreg/_0573_ ), .Z(\myreg/_3023_ ) );
BUF_X1 \myreg/_6562_ ( .A(\myreg/_0574_ ), .Z(\myreg/_3024_ ) );
BUF_X1 \myreg/_6563_ ( .A(\myreg/_0575_ ), .Z(\myreg/_3025_ ) );
BUF_X1 \myreg/_6564_ ( .A(\myreg/_0576_ ), .Z(\myreg/_3026_ ) );
BUF_X1 \myreg/_6565_ ( .A(\myreg/_0577_ ), .Z(\myreg/_3027_ ) );
BUF_X1 \myreg/_6566_ ( .A(\myreg/_0578_ ), .Z(\myreg/_3028_ ) );
BUF_X1 \myreg/_6567_ ( .A(\myreg/_0579_ ), .Z(\myreg/_3029_ ) );
BUF_X1 \myreg/_6568_ ( .A(\myreg/_0580_ ), .Z(\myreg/_3030_ ) );
BUF_X1 \myreg/_6569_ ( .A(\myreg/_0581_ ), .Z(\myreg/_3031_ ) );
BUF_X1 \myreg/_6570_ ( .A(\myreg/_0582_ ), .Z(\myreg/_3032_ ) );
BUF_X1 \myreg/_6571_ ( .A(\myreg/_0583_ ), .Z(\myreg/_3033_ ) );
BUF_X1 \myreg/_6572_ ( .A(\myreg/_0584_ ), .Z(\myreg/_3034_ ) );
BUF_X1 \myreg/_6573_ ( .A(\myreg/_0585_ ), .Z(\myreg/_3035_ ) );
BUF_X1 \myreg/_6574_ ( .A(\myreg/_0586_ ), .Z(\myreg/_3036_ ) );
BUF_X1 \myreg/_6575_ ( .A(\myreg/_0587_ ), .Z(\myreg/_3037_ ) );
BUF_X1 \myreg/_6576_ ( .A(\myreg/_0588_ ), .Z(\myreg/_3038_ ) );
BUF_X1 \myreg/_6577_ ( .A(\myreg/_0589_ ), .Z(\myreg/_3039_ ) );
BUF_X1 \myreg/_6578_ ( .A(\myreg/_0590_ ), .Z(\myreg/_3040_ ) );
BUF_X1 \myreg/_6579_ ( .A(\myreg/_0591_ ), .Z(\myreg/_3041_ ) );
BUF_X1 \myreg/_6580_ ( .A(\myreg/_0592_ ), .Z(\myreg/_3042_ ) );
BUF_X1 \myreg/_6581_ ( .A(\myreg/_0593_ ), .Z(\myreg/_3043_ ) );
BUF_X1 \myreg/_6582_ ( .A(\myreg/_0594_ ), .Z(\myreg/_3044_ ) );
BUF_X1 \myreg/_6583_ ( .A(\myreg/_0595_ ), .Z(\myreg/_3045_ ) );
BUF_X1 \myreg/_6584_ ( .A(\myreg/_0596_ ), .Z(\myreg/_3046_ ) );
BUF_X1 \myreg/_6585_ ( .A(\myreg/_0597_ ), .Z(\myreg/_3047_ ) );
BUF_X1 \myreg/_6586_ ( .A(\myreg/_0598_ ), .Z(\myreg/_3048_ ) );
BUF_X1 \myreg/_6587_ ( .A(\myreg/_0599_ ), .Z(\myreg/_3049_ ) );
BUF_X1 \myreg/_6588_ ( .A(\myreg/_0600_ ), .Z(\myreg/_3050_ ) );
BUF_X1 \myreg/_6589_ ( .A(\myreg/_0601_ ), .Z(\myreg/_3051_ ) );
BUF_X1 \myreg/_6590_ ( .A(\myreg/_0602_ ), .Z(\myreg/_3052_ ) );
BUF_X1 \myreg/_6591_ ( .A(\myreg/_0603_ ), .Z(\myreg/_3053_ ) );
BUF_X1 \myreg/_6592_ ( .A(\myreg/_0604_ ), .Z(\myreg/_3054_ ) );
BUF_X1 \myreg/_6593_ ( .A(\myreg/_0605_ ), .Z(\myreg/_3055_ ) );
BUF_X1 \myreg/_6594_ ( .A(\myreg/_0606_ ), .Z(\myreg/_3056_ ) );
BUF_X1 \myreg/_6595_ ( .A(\myreg/_0607_ ), .Z(\myreg/_3057_ ) );
BUF_X1 \myreg/_6596_ ( .A(\myreg/_0608_ ), .Z(\myreg/_3058_ ) );
BUF_X1 \myreg/_6597_ ( .A(\myreg/_0609_ ), .Z(\myreg/_3059_ ) );
BUF_X1 \myreg/_6598_ ( .A(\myreg/_0610_ ), .Z(\myreg/_3060_ ) );
BUF_X1 \myreg/_6599_ ( .A(\myreg/_0611_ ), .Z(\myreg/_3061_ ) );
BUF_X1 \myreg/_6600_ ( .A(\myreg/_0612_ ), .Z(\myreg/_3062_ ) );
BUF_X1 \myreg/_6601_ ( .A(\myreg/_0613_ ), .Z(\myreg/_3063_ ) );
BUF_X1 \myreg/_6602_ ( .A(\myreg/_0614_ ), .Z(\myreg/_3064_ ) );
BUF_X1 \myreg/_6603_ ( .A(\myreg/_0615_ ), .Z(\myreg/_3065_ ) );
BUF_X1 \myreg/_6604_ ( .A(\myreg/_0616_ ), .Z(\myreg/_3066_ ) );
BUF_X1 \myreg/_6605_ ( .A(\myreg/_0617_ ), .Z(\myreg/_3067_ ) );
BUF_X1 \myreg/_6606_ ( .A(\myreg/_0618_ ), .Z(\myreg/_3068_ ) );
BUF_X1 \myreg/_6607_ ( .A(\myreg/_0619_ ), .Z(\myreg/_3069_ ) );
BUF_X1 \myreg/_6608_ ( .A(\myreg/_0620_ ), .Z(\myreg/_3070_ ) );
BUF_X1 \myreg/_6609_ ( .A(\myreg/_0621_ ), .Z(\myreg/_3071_ ) );
BUF_X1 \myreg/_6610_ ( .A(\myreg/_0622_ ), .Z(\myreg/_3072_ ) );
BUF_X1 \myreg/_6611_ ( .A(\myreg/_0623_ ), .Z(\myreg/_3073_ ) );
BUF_X1 \myreg/_6612_ ( .A(\myreg/_0624_ ), .Z(\myreg/_3074_ ) );
BUF_X1 \myreg/_6613_ ( .A(\myreg/_0625_ ), .Z(\myreg/_3075_ ) );
BUF_X1 \myreg/_6614_ ( .A(\myreg/_0626_ ), .Z(\myreg/_3076_ ) );
BUF_X1 \myreg/_6615_ ( .A(\myreg/_0627_ ), .Z(\myreg/_3077_ ) );
BUF_X1 \myreg/_6616_ ( .A(\myreg/_0628_ ), .Z(\myreg/_3078_ ) );
BUF_X1 \myreg/_6617_ ( .A(\myreg/_0629_ ), .Z(\myreg/_3079_ ) );
BUF_X1 \myreg/_6618_ ( .A(\myreg/_0630_ ), .Z(\myreg/_3080_ ) );
BUF_X1 \myreg/_6619_ ( .A(\myreg/_0631_ ), .Z(\myreg/_3081_ ) );
BUF_X1 \myreg/_6620_ ( .A(\myreg/_0632_ ), .Z(\myreg/_3082_ ) );
BUF_X1 \myreg/_6621_ ( .A(\myreg/_0633_ ), .Z(\myreg/_3083_ ) );
BUF_X1 \myreg/_6622_ ( .A(\myreg/_0634_ ), .Z(\myreg/_3084_ ) );
BUF_X1 \myreg/_6623_ ( .A(\myreg/_0635_ ), .Z(\myreg/_3085_ ) );
BUF_X1 \myreg/_6624_ ( .A(\myreg/_0636_ ), .Z(\myreg/_3086_ ) );
BUF_X1 \myreg/_6625_ ( .A(\myreg/_0637_ ), .Z(\myreg/_3087_ ) );
BUF_X1 \myreg/_6626_ ( .A(\myreg/_0638_ ), .Z(\myreg/_3088_ ) );
BUF_X1 \myreg/_6627_ ( .A(\myreg/_0639_ ), .Z(\myreg/_3089_ ) );
BUF_X1 \myreg/_6628_ ( .A(\myreg/_0640_ ), .Z(\myreg/_3090_ ) );
BUF_X1 \myreg/_6629_ ( .A(\myreg/_0641_ ), .Z(\myreg/_3091_ ) );
BUF_X1 \myreg/_6630_ ( .A(\myreg/_0642_ ), .Z(\myreg/_3092_ ) );
BUF_X1 \myreg/_6631_ ( .A(\myreg/_0643_ ), .Z(\myreg/_3093_ ) );
BUF_X1 \myreg/_6632_ ( .A(\myreg/_0644_ ), .Z(\myreg/_3094_ ) );
BUF_X1 \myreg/_6633_ ( .A(\myreg/_0645_ ), .Z(\myreg/_3095_ ) );
BUF_X1 \myreg/_6634_ ( .A(\myreg/_0646_ ), .Z(\myreg/_3096_ ) );
BUF_X1 \myreg/_6635_ ( .A(\myreg/_0647_ ), .Z(\myreg/_3097_ ) );
BUF_X1 \myreg/_6636_ ( .A(\myreg/_0648_ ), .Z(\myreg/_3098_ ) );
BUF_X1 \myreg/_6637_ ( .A(\myreg/_0649_ ), .Z(\myreg/_3099_ ) );
BUF_X1 \myreg/_6638_ ( .A(\myreg/_0650_ ), .Z(\myreg/_3100_ ) );
BUF_X1 \myreg/_6639_ ( .A(\myreg/_0651_ ), .Z(\myreg/_3101_ ) );
BUF_X1 \myreg/_6640_ ( .A(\myreg/_0652_ ), .Z(\myreg/_3102_ ) );
BUF_X1 \myreg/_6641_ ( .A(\myreg/_0653_ ), .Z(\myreg/_3103_ ) );
BUF_X1 \myreg/_6642_ ( .A(\myreg/_0654_ ), .Z(\myreg/_3104_ ) );
BUF_X1 \myreg/_6643_ ( .A(\myreg/_0655_ ), .Z(\myreg/_3105_ ) );
BUF_X1 \myreg/_6644_ ( .A(\myreg/_0656_ ), .Z(\myreg/_3106_ ) );
BUF_X1 \myreg/_6645_ ( .A(\myreg/_0657_ ), .Z(\myreg/_3107_ ) );
BUF_X1 \myreg/_6646_ ( .A(\myreg/_0658_ ), .Z(\myreg/_3108_ ) );
BUF_X1 \myreg/_6647_ ( .A(\myreg/_0659_ ), .Z(\myreg/_3109_ ) );
BUF_X1 \myreg/_6648_ ( .A(\myreg/_0660_ ), .Z(\myreg/_3110_ ) );
BUF_X1 \myreg/_6649_ ( .A(\myreg/_0661_ ), .Z(\myreg/_3111_ ) );
BUF_X1 \myreg/_6650_ ( .A(\myreg/_0662_ ), .Z(\myreg/_3112_ ) );
BUF_X1 \myreg/_6651_ ( .A(\myreg/_0663_ ), .Z(\myreg/_3113_ ) );
BUF_X1 \myreg/_6652_ ( .A(\myreg/_0664_ ), .Z(\myreg/_3114_ ) );
BUF_X1 \myreg/_6653_ ( .A(\myreg/_0665_ ), .Z(\myreg/_3115_ ) );
BUF_X1 \myreg/_6654_ ( .A(\myreg/_0666_ ), .Z(\myreg/_3116_ ) );
BUF_X1 \myreg/_6655_ ( .A(\myreg/_0667_ ), .Z(\myreg/_3117_ ) );
BUF_X1 \myreg/_6656_ ( .A(\myreg/_0668_ ), .Z(\myreg/_3118_ ) );
BUF_X1 \myreg/_6657_ ( .A(\myreg/_0669_ ), .Z(\myreg/_3119_ ) );
BUF_X1 \myreg/_6658_ ( .A(\myreg/_0670_ ), .Z(\myreg/_3120_ ) );
BUF_X1 \myreg/_6659_ ( .A(\myreg/_0671_ ), .Z(\myreg/_3121_ ) );
BUF_X1 \myreg/_6660_ ( .A(\myreg/_0672_ ), .Z(\myreg/_3122_ ) );
BUF_X1 \myreg/_6661_ ( .A(\myreg/_0673_ ), .Z(\myreg/_3123_ ) );
BUF_X1 \myreg/_6662_ ( .A(\myreg/_0674_ ), .Z(\myreg/_3124_ ) );
BUF_X1 \myreg/_6663_ ( .A(\myreg/_0675_ ), .Z(\myreg/_3125_ ) );
BUF_X1 \myreg/_6664_ ( .A(\myreg/_0676_ ), .Z(\myreg/_3126_ ) );
BUF_X1 \myreg/_6665_ ( .A(\myreg/_0677_ ), .Z(\myreg/_3127_ ) );
BUF_X1 \myreg/_6666_ ( .A(\myreg/_0678_ ), .Z(\myreg/_3128_ ) );
BUF_X1 \myreg/_6667_ ( .A(\myreg/_0679_ ), .Z(\myreg/_3129_ ) );
BUF_X1 \myreg/_6668_ ( .A(\myreg/_0680_ ), .Z(\myreg/_3130_ ) );
BUF_X1 \myreg/_6669_ ( .A(\myreg/_0681_ ), .Z(\myreg/_3131_ ) );
BUF_X1 \myreg/_6670_ ( .A(\myreg/_0682_ ), .Z(\myreg/_3132_ ) );
BUF_X1 \myreg/_6671_ ( .A(\myreg/_0683_ ), .Z(\myreg/_3133_ ) );
BUF_X1 \myreg/_6672_ ( .A(\myreg/_0684_ ), .Z(\myreg/_3134_ ) );
BUF_X1 \myreg/_6673_ ( .A(\myreg/_0685_ ), .Z(\myreg/_3135_ ) );
BUF_X1 \myreg/_6674_ ( .A(\myreg/_0686_ ), .Z(\myreg/_3136_ ) );
BUF_X1 \myreg/_6675_ ( .A(\myreg/_0687_ ), .Z(\myreg/_3137_ ) );
BUF_X1 \myreg/_6676_ ( .A(\myreg/_0688_ ), .Z(\myreg/_3138_ ) );
BUF_X1 \myreg/_6677_ ( .A(\myreg/_0689_ ), .Z(\myreg/_3139_ ) );
BUF_X1 \myreg/_6678_ ( .A(\myreg/_0690_ ), .Z(\myreg/_3140_ ) );
BUF_X1 \myreg/_6679_ ( .A(\myreg/_0691_ ), .Z(\myreg/_3141_ ) );
BUF_X1 \myreg/_6680_ ( .A(\myreg/_0692_ ), .Z(\myreg/_3142_ ) );
BUF_X1 \myreg/_6681_ ( .A(\myreg/_0693_ ), .Z(\myreg/_3143_ ) );
BUF_X1 \myreg/_6682_ ( .A(\myreg/_0694_ ), .Z(\myreg/_3144_ ) );
BUF_X1 \myreg/_6683_ ( .A(\myreg/_0695_ ), .Z(\myreg/_3145_ ) );
BUF_X1 \myreg/_6684_ ( .A(\myreg/_0696_ ), .Z(\myreg/_3146_ ) );
BUF_X1 \myreg/_6685_ ( .A(\myreg/_0697_ ), .Z(\myreg/_3147_ ) );
BUF_X1 \myreg/_6686_ ( .A(\myreg/_0698_ ), .Z(\myreg/_3148_ ) );
BUF_X1 \myreg/_6687_ ( .A(\myreg/_0699_ ), .Z(\myreg/_3149_ ) );
BUF_X1 \myreg/_6688_ ( .A(\myreg/_0700_ ), .Z(\myreg/_3150_ ) );
BUF_X1 \myreg/_6689_ ( .A(\myreg/_0701_ ), .Z(\myreg/_3151_ ) );
BUF_X1 \myreg/_6690_ ( .A(\myreg/_0702_ ), .Z(\myreg/_3152_ ) );
BUF_X1 \myreg/_6691_ ( .A(\myreg/_0703_ ), .Z(\myreg/_3153_ ) );
BUF_X1 \myreg/_6692_ ( .A(\myreg/_0704_ ), .Z(\myreg/_3154_ ) );
BUF_X1 \myreg/_6693_ ( .A(\myreg/_0705_ ), .Z(\myreg/_3155_ ) );
BUF_X1 \myreg/_6694_ ( .A(\myreg/_0706_ ), .Z(\myreg/_3156_ ) );
BUF_X1 \myreg/_6695_ ( .A(\myreg/_0707_ ), .Z(\myreg/_3157_ ) );
BUF_X1 \myreg/_6696_ ( .A(\myreg/_0708_ ), .Z(\myreg/_3158_ ) );
BUF_X1 \myreg/_6697_ ( .A(\myreg/_0709_ ), .Z(\myreg/_3159_ ) );
BUF_X1 \myreg/_6698_ ( .A(\myreg/_0710_ ), .Z(\myreg/_3160_ ) );
BUF_X1 \myreg/_6699_ ( .A(\myreg/_0711_ ), .Z(\myreg/_3161_ ) );
BUF_X1 \myreg/_6700_ ( .A(\myreg/_0712_ ), .Z(\myreg/_3162_ ) );
BUF_X1 \myreg/_6701_ ( .A(\myreg/_0713_ ), .Z(\myreg/_3163_ ) );
BUF_X1 \myreg/_6702_ ( .A(\myreg/_0714_ ), .Z(\myreg/_3164_ ) );
BUF_X1 \myreg/_6703_ ( .A(\myreg/_0715_ ), .Z(\myreg/_3165_ ) );
BUF_X1 \myreg/_6704_ ( .A(\myreg/_0716_ ), .Z(\myreg/_3166_ ) );
BUF_X1 \myreg/_6705_ ( .A(\myreg/_0717_ ), .Z(\myreg/_3167_ ) );
BUF_X1 \myreg/_6706_ ( .A(\myreg/_0718_ ), .Z(\myreg/_3168_ ) );
BUF_X1 \myreg/_6707_ ( .A(\myreg/_0719_ ), .Z(\myreg/_3169_ ) );
BUF_X1 \myreg/_6708_ ( .A(\myreg/_0720_ ), .Z(\myreg/_3170_ ) );
BUF_X1 \myreg/_6709_ ( .A(\myreg/_0721_ ), .Z(\myreg/_3171_ ) );
BUF_X1 \myreg/_6710_ ( .A(\myreg/_0722_ ), .Z(\myreg/_3172_ ) );
BUF_X1 \myreg/_6711_ ( .A(\myreg/_0723_ ), .Z(\myreg/_3173_ ) );
BUF_X1 \myreg/_6712_ ( .A(\myreg/_0724_ ), .Z(\myreg/_3174_ ) );
BUF_X1 \myreg/_6713_ ( .A(\myreg/_0725_ ), .Z(\myreg/_3175_ ) );
BUF_X1 \myreg/_6714_ ( .A(\myreg/_0726_ ), .Z(\myreg/_3176_ ) );
BUF_X1 \myreg/_6715_ ( .A(\myreg/_0727_ ), .Z(\myreg/_3177_ ) );
BUF_X1 \myreg/_6716_ ( .A(\myreg/_0728_ ), .Z(\myreg/_3178_ ) );
BUF_X1 \myreg/_6717_ ( .A(\myreg/_0729_ ), .Z(\myreg/_3179_ ) );
BUF_X1 \myreg/_6718_ ( .A(\myreg/_0730_ ), .Z(\myreg/_3180_ ) );
BUF_X1 \myreg/_6719_ ( .A(\myreg/_0731_ ), .Z(\myreg/_3181_ ) );
BUF_X1 \myreg/_6720_ ( .A(\myreg/_0732_ ), .Z(\myreg/_3182_ ) );
BUF_X1 \myreg/_6721_ ( .A(\myreg/_0733_ ), .Z(\myreg/_3183_ ) );
BUF_X1 \myreg/_6722_ ( .A(\myreg/_0734_ ), .Z(\myreg/_3184_ ) );
BUF_X1 \myreg/_6723_ ( .A(\myreg/_0735_ ), .Z(\myreg/_3185_ ) );
BUF_X1 \myreg/_6724_ ( .A(\myreg/_0736_ ), .Z(\myreg/_3186_ ) );
BUF_X1 \myreg/_6725_ ( .A(\myreg/_0737_ ), .Z(\myreg/_3187_ ) );
BUF_X1 \myreg/_6726_ ( .A(\myreg/_0738_ ), .Z(\myreg/_3188_ ) );
BUF_X1 \myreg/_6727_ ( .A(\myreg/_0739_ ), .Z(\myreg/_3189_ ) );
BUF_X1 \myreg/_6728_ ( .A(\myreg/_0740_ ), .Z(\myreg/_3190_ ) );
BUF_X1 \myreg/_6729_ ( .A(\myreg/_0741_ ), .Z(\myreg/_3191_ ) );
BUF_X1 \myreg/_6730_ ( .A(\myreg/_0742_ ), .Z(\myreg/_3192_ ) );
BUF_X1 \myreg/_6731_ ( .A(\myreg/_0743_ ), .Z(\myreg/_3193_ ) );
BUF_X1 \myreg/_6732_ ( .A(\myreg/_0744_ ), .Z(\myreg/_3194_ ) );
BUF_X1 \myreg/_6733_ ( .A(\myreg/_0745_ ), .Z(\myreg/_3195_ ) );
BUF_X1 \myreg/_6734_ ( .A(\myreg/_0746_ ), .Z(\myreg/_3196_ ) );
BUF_X1 \myreg/_6735_ ( .A(\myreg/_0747_ ), .Z(\myreg/_3197_ ) );
BUF_X1 \myreg/_6736_ ( .A(\myreg/_0748_ ), .Z(\myreg/_3198_ ) );
BUF_X1 \myreg/_6737_ ( .A(\myreg/_0749_ ), .Z(\myreg/_3199_ ) );
BUF_X1 \myreg/_6738_ ( .A(\myreg/_0750_ ), .Z(\myreg/_3200_ ) );
BUF_X1 \myreg/_6739_ ( .A(\myreg/_0751_ ), .Z(\myreg/_3201_ ) );
BUF_X1 \myreg/_6740_ ( .A(\myreg/_0752_ ), .Z(\myreg/_3202_ ) );
BUF_X1 \myreg/_6741_ ( .A(\myreg/_0753_ ), .Z(\myreg/_3203_ ) );
BUF_X1 \myreg/_6742_ ( .A(\myreg/_0754_ ), .Z(\myreg/_3204_ ) );
BUF_X1 \myreg/_6743_ ( .A(\myreg/_0755_ ), .Z(\myreg/_3205_ ) );
BUF_X1 \myreg/_6744_ ( .A(\myreg/_0756_ ), .Z(\myreg/_3206_ ) );
BUF_X1 \myreg/_6745_ ( .A(\myreg/_0757_ ), .Z(\myreg/_3207_ ) );
BUF_X1 \myreg/_6746_ ( .A(\myreg/_0758_ ), .Z(\myreg/_3208_ ) );
BUF_X1 \myreg/_6747_ ( .A(\myreg/_0759_ ), .Z(\myreg/_3209_ ) );
BUF_X1 \myreg/_6748_ ( .A(\myreg/_0760_ ), .Z(\myreg/_3210_ ) );
BUF_X1 \myreg/_6749_ ( .A(\myreg/_0761_ ), .Z(\myreg/_3211_ ) );
BUF_X1 \myreg/_6750_ ( .A(\myreg/_0762_ ), .Z(\myreg/_3212_ ) );
BUF_X1 \myreg/_6751_ ( .A(\myreg/_0763_ ), .Z(\myreg/_3213_ ) );
BUF_X1 \myreg/_6752_ ( .A(\myreg/_0764_ ), .Z(\myreg/_3214_ ) );
BUF_X1 \myreg/_6753_ ( .A(\myreg/_0765_ ), .Z(\myreg/_3215_ ) );
BUF_X1 \myreg/_6754_ ( .A(\myreg/_0766_ ), .Z(\myreg/_3216_ ) );
BUF_X1 \myreg/_6755_ ( .A(\myreg/_0767_ ), .Z(\myreg/_3217_ ) );
BUF_X1 \myreg/_6756_ ( .A(\myreg/_0768_ ), .Z(\myreg/_3218_ ) );
BUF_X1 \myreg/_6757_ ( .A(\myreg/_0769_ ), .Z(\myreg/_3219_ ) );
BUF_X1 \myreg/_6758_ ( .A(\myreg/_0770_ ), .Z(\myreg/_3220_ ) );
BUF_X1 \myreg/_6759_ ( .A(\myreg/_0771_ ), .Z(\myreg/_3221_ ) );
BUF_X1 \myreg/_6760_ ( .A(\myreg/_0772_ ), .Z(\myreg/_3222_ ) );
BUF_X1 \myreg/_6761_ ( .A(\myreg/_0773_ ), .Z(\myreg/_3223_ ) );
BUF_X1 \myreg/_6762_ ( .A(\myreg/_0774_ ), .Z(\myreg/_3224_ ) );
BUF_X1 \myreg/_6763_ ( .A(\myreg/_0775_ ), .Z(\myreg/_3225_ ) );
BUF_X1 \myreg/_6764_ ( .A(\myreg/_0776_ ), .Z(\myreg/_3226_ ) );
BUF_X1 \myreg/_6765_ ( .A(\myreg/_0777_ ), .Z(\myreg/_3227_ ) );
BUF_X1 \myreg/_6766_ ( .A(\myreg/_0778_ ), .Z(\myreg/_3228_ ) );
BUF_X1 \myreg/_6767_ ( .A(\myreg/_0779_ ), .Z(\myreg/_3229_ ) );
BUF_X1 \myreg/_6768_ ( .A(\myreg/_0780_ ), .Z(\myreg/_3230_ ) );
BUF_X1 \myreg/_6769_ ( .A(\myreg/_0781_ ), .Z(\myreg/_3231_ ) );
BUF_X1 \myreg/_6770_ ( .A(\myreg/_0782_ ), .Z(\myreg/_3232_ ) );
BUF_X1 \myreg/_6771_ ( .A(\myreg/_0783_ ), .Z(\myreg/_3233_ ) );
BUF_X1 \myreg/_6772_ ( .A(\myreg/_0784_ ), .Z(\myreg/_3234_ ) );
BUF_X1 \myreg/_6773_ ( .A(\myreg/_0785_ ), .Z(\myreg/_3235_ ) );
BUF_X1 \myreg/_6774_ ( .A(\myreg/_0786_ ), .Z(\myreg/_3236_ ) );
BUF_X1 \myreg/_6775_ ( .A(\myreg/_0787_ ), .Z(\myreg/_3237_ ) );
BUF_X1 \myreg/_6776_ ( .A(\myreg/_0788_ ), .Z(\myreg/_3238_ ) );
BUF_X1 \myreg/_6777_ ( .A(\myreg/_0789_ ), .Z(\myreg/_3239_ ) );
BUF_X1 \myreg/_6778_ ( .A(\myreg/_0790_ ), .Z(\myreg/_3240_ ) );
BUF_X1 \myreg/_6779_ ( .A(\myreg/_0791_ ), .Z(\myreg/_3241_ ) );
BUF_X1 \myreg/_6780_ ( .A(\myreg/_0792_ ), .Z(\myreg/_3242_ ) );
BUF_X1 \myreg/_6781_ ( .A(\myreg/_0793_ ), .Z(\myreg/_3243_ ) );
BUF_X1 \myreg/_6782_ ( .A(\myreg/_0794_ ), .Z(\myreg/_3244_ ) );
BUF_X1 \myreg/_6783_ ( .A(\myreg/_0795_ ), .Z(\myreg/_3245_ ) );
BUF_X1 \myreg/_6784_ ( .A(\myreg/_0796_ ), .Z(\myreg/_3246_ ) );
BUF_X1 \myreg/_6785_ ( .A(\myreg/_0797_ ), .Z(\myreg/_3247_ ) );
BUF_X1 \myreg/_6786_ ( .A(\myreg/_0798_ ), .Z(\myreg/_3248_ ) );
BUF_X1 \myreg/_6787_ ( .A(\myreg/_0799_ ), .Z(\myreg/_3249_ ) );
BUF_X1 \myreg/_6788_ ( .A(\myreg/_0800_ ), .Z(\myreg/_3250_ ) );
BUF_X1 \myreg/_6789_ ( .A(\myreg/_0801_ ), .Z(\myreg/_3251_ ) );
BUF_X1 \myreg/_6790_ ( .A(\myreg/_0802_ ), .Z(\myreg/_3252_ ) );
BUF_X1 \myreg/_6791_ ( .A(\myreg/_0803_ ), .Z(\myreg/_3253_ ) );
BUF_X1 \myreg/_6792_ ( .A(\myreg/_0804_ ), .Z(\myreg/_3254_ ) );
BUF_X1 \myreg/_6793_ ( .A(\myreg/_0805_ ), .Z(\myreg/_3255_ ) );
BUF_X1 \myreg/_6794_ ( .A(\myreg/_0806_ ), .Z(\myreg/_3256_ ) );
BUF_X1 \myreg/_6795_ ( .A(\myreg/_0807_ ), .Z(\myreg/_3257_ ) );
BUF_X1 \myreg/_6796_ ( .A(\myreg/_0808_ ), .Z(\myreg/_3258_ ) );
BUF_X1 \myreg/_6797_ ( .A(\myreg/_0809_ ), .Z(\myreg/_3259_ ) );
BUF_X1 \myreg/_6798_ ( .A(\myreg/_0810_ ), .Z(\myreg/_3260_ ) );
BUF_X1 \myreg/_6799_ ( .A(\myreg/_0811_ ), .Z(\myreg/_3261_ ) );
BUF_X1 \myreg/_6800_ ( .A(\myreg/_0812_ ), .Z(\myreg/_3262_ ) );
BUF_X1 \myreg/_6801_ ( .A(\myreg/_0813_ ), .Z(\myreg/_3263_ ) );
BUF_X1 \myreg/_6802_ ( .A(\myreg/_0814_ ), .Z(\myreg/_3264_ ) );
BUF_X1 \myreg/_6803_ ( .A(\myreg/_0815_ ), .Z(\myreg/_3265_ ) );
BUF_X1 \myreg/_6804_ ( .A(\myreg/_0816_ ), .Z(\myreg/_3266_ ) );
BUF_X1 \myreg/_6805_ ( .A(\myreg/_0817_ ), .Z(\myreg/_3267_ ) );
BUF_X1 \myreg/_6806_ ( .A(\myreg/_0818_ ), .Z(\myreg/_3268_ ) );
BUF_X1 \myreg/_6807_ ( .A(\myreg/_0819_ ), .Z(\myreg/_3269_ ) );
BUF_X1 \myreg/_6808_ ( .A(\myreg/_0820_ ), .Z(\myreg/_3270_ ) );
BUF_X1 \myreg/_6809_ ( .A(\myreg/_0821_ ), .Z(\myreg/_3271_ ) );
BUF_X1 \myreg/_6810_ ( .A(\myreg/_0822_ ), .Z(\myreg/_3272_ ) );
BUF_X1 \myreg/_6811_ ( .A(\myreg/_0823_ ), .Z(\myreg/_3273_ ) );
BUF_X1 \myreg/_6812_ ( .A(\myreg/_0824_ ), .Z(\myreg/_3274_ ) );
BUF_X1 \myreg/_6813_ ( .A(\myreg/_0825_ ), .Z(\myreg/_3275_ ) );
BUF_X1 \myreg/_6814_ ( .A(\myreg/_0826_ ), .Z(\myreg/_3276_ ) );
BUF_X1 \myreg/_6815_ ( .A(\myreg/_0827_ ), .Z(\myreg/_3277_ ) );
BUF_X1 \myreg/_6816_ ( .A(\myreg/_0828_ ), .Z(\myreg/_3278_ ) );
BUF_X1 \myreg/_6817_ ( .A(\myreg/_0829_ ), .Z(\myreg/_3279_ ) );
BUF_X1 \myreg/_6818_ ( .A(\myreg/_0830_ ), .Z(\myreg/_3280_ ) );
BUF_X1 \myreg/_6819_ ( .A(\myreg/_0831_ ), .Z(\myreg/_3281_ ) );
BUF_X1 \myreg/_6820_ ( .A(\myreg/_0832_ ), .Z(\myreg/_3282_ ) );
BUF_X1 \myreg/_6821_ ( .A(\myreg/_0833_ ), .Z(\myreg/_3283_ ) );
BUF_X1 \myreg/_6822_ ( .A(\myreg/_0834_ ), .Z(\myreg/_3284_ ) );
BUF_X1 \myreg/_6823_ ( .A(\myreg/_0835_ ), .Z(\myreg/_3285_ ) );
BUF_X1 \myreg/_6824_ ( .A(\myreg/_0836_ ), .Z(\myreg/_3286_ ) );
BUF_X1 \myreg/_6825_ ( .A(\myreg/_0837_ ), .Z(\myreg/_3287_ ) );
BUF_X1 \myreg/_6826_ ( .A(\myreg/_0838_ ), .Z(\myreg/_3288_ ) );
BUF_X1 \myreg/_6827_ ( .A(\myreg/_0839_ ), .Z(\myreg/_3289_ ) );
BUF_X1 \myreg/_6828_ ( .A(\myreg/_0840_ ), .Z(\myreg/_3290_ ) );
BUF_X1 \myreg/_6829_ ( .A(\myreg/_0841_ ), .Z(\myreg/_3291_ ) );
BUF_X1 \myreg/_6830_ ( .A(\myreg/_0842_ ), .Z(\myreg/_3292_ ) );
BUF_X1 \myreg/_6831_ ( .A(\myreg/_0843_ ), .Z(\myreg/_3293_ ) );
BUF_X1 \myreg/_6832_ ( .A(\myreg/_0844_ ), .Z(\myreg/_3294_ ) );
BUF_X1 \myreg/_6833_ ( .A(\myreg/_0845_ ), .Z(\myreg/_3295_ ) );
BUF_X1 \myreg/_6834_ ( .A(\myreg/_0846_ ), .Z(\myreg/_3296_ ) );
BUF_X1 \myreg/_6835_ ( .A(\myreg/_0847_ ), .Z(\myreg/_3297_ ) );
BUF_X1 \myreg/_6836_ ( .A(\myreg/_0848_ ), .Z(\myreg/_3298_ ) );
BUF_X1 \myreg/_6837_ ( .A(\myreg/_0849_ ), .Z(\myreg/_3299_ ) );
BUF_X1 \myreg/_6838_ ( .A(\myreg/_0850_ ), .Z(\myreg/_3300_ ) );
BUF_X1 \myreg/_6839_ ( .A(\myreg/_0851_ ), .Z(\myreg/_3301_ ) );
BUF_X1 \myreg/_6840_ ( .A(\myreg/_0852_ ), .Z(\myreg/_3302_ ) );
BUF_X1 \myreg/_6841_ ( .A(\myreg/_0853_ ), .Z(\myreg/_3303_ ) );
BUF_X1 \myreg/_6842_ ( .A(\myreg/_0854_ ), .Z(\myreg/_3304_ ) );
BUF_X1 \myreg/_6843_ ( .A(\myreg/_0855_ ), .Z(\myreg/_3305_ ) );
BUF_X1 \myreg/_6844_ ( .A(\myreg/_0856_ ), .Z(\myreg/_3306_ ) );
BUF_X1 \myreg/_6845_ ( .A(\myreg/_0857_ ), .Z(\myreg/_3307_ ) );
BUF_X1 \myreg/_6846_ ( .A(\myreg/_0858_ ), .Z(\myreg/_3308_ ) );
BUF_X1 \myreg/_6847_ ( .A(\myreg/_0859_ ), .Z(\myreg/_3309_ ) );
BUF_X1 \myreg/_6848_ ( .A(\myreg/_0860_ ), .Z(\myreg/_3310_ ) );
BUF_X1 \myreg/_6849_ ( .A(\myreg/_0861_ ), .Z(\myreg/_3311_ ) );
BUF_X1 \myreg/_6850_ ( .A(\myreg/_0862_ ), .Z(\myreg/_3312_ ) );
BUF_X1 \myreg/_6851_ ( .A(\myreg/_0863_ ), .Z(\myreg/_3313_ ) );
BUF_X1 \myreg/_6852_ ( .A(\myreg/_0864_ ), .Z(\myreg/_3314_ ) );
BUF_X1 \myreg/_6853_ ( .A(\myreg/_0865_ ), .Z(\myreg/_3315_ ) );
BUF_X1 \myreg/_6854_ ( .A(\myreg/_0866_ ), .Z(\myreg/_3316_ ) );
BUF_X1 \myreg/_6855_ ( .A(\myreg/_0867_ ), .Z(\myreg/_3317_ ) );
BUF_X1 \myreg/_6856_ ( .A(\myreg/_0868_ ), .Z(\myreg/_3318_ ) );
BUF_X1 \myreg/_6857_ ( .A(\myreg/_0869_ ), .Z(\myreg/_3319_ ) );
BUF_X1 \myreg/_6858_ ( .A(\myreg/_0870_ ), .Z(\myreg/_3320_ ) );
BUF_X1 \myreg/_6859_ ( .A(\myreg/_0871_ ), .Z(\myreg/_3321_ ) );
BUF_X1 \myreg/_6860_ ( .A(\myreg/_0872_ ), .Z(\myreg/_3322_ ) );
BUF_X1 \myreg/_6861_ ( .A(\myreg/_0873_ ), .Z(\myreg/_3323_ ) );
BUF_X1 \myreg/_6862_ ( .A(\myreg/_0874_ ), .Z(\myreg/_3324_ ) );
BUF_X1 \myreg/_6863_ ( .A(\myreg/_0875_ ), .Z(\myreg/_3325_ ) );
BUF_X1 \myreg/_6864_ ( .A(\myreg/_0876_ ), .Z(\myreg/_3326_ ) );
BUF_X1 \myreg/_6865_ ( .A(\myreg/_0877_ ), .Z(\myreg/_3327_ ) );
BUF_X1 \myreg/_6866_ ( .A(\myreg/_0878_ ), .Z(\myreg/_3328_ ) );
BUF_X1 \myreg/_6867_ ( .A(\myreg/_0879_ ), .Z(\myreg/_3329_ ) );
BUF_X1 \myreg/_6868_ ( .A(\myreg/_0880_ ), .Z(\myreg/_3330_ ) );
BUF_X1 \myreg/_6869_ ( .A(\myreg/_0881_ ), .Z(\myreg/_3331_ ) );
BUF_X1 \myreg/_6870_ ( .A(\myreg/_0882_ ), .Z(\myreg/_3332_ ) );
BUF_X1 \myreg/_6871_ ( .A(\myreg/_0883_ ), .Z(\myreg/_3333_ ) );
BUF_X1 \myreg/_6872_ ( .A(\myreg/_0884_ ), .Z(\myreg/_3334_ ) );
BUF_X1 \myreg/_6873_ ( .A(\myreg/_0885_ ), .Z(\myreg/_3335_ ) );
BUF_X1 \myreg/_6874_ ( .A(\myreg/_0886_ ), .Z(\myreg/_3336_ ) );
BUF_X1 \myreg/_6875_ ( .A(\myreg/_0887_ ), .Z(\myreg/_3337_ ) );
BUF_X1 \myreg/_6876_ ( .A(\myreg/_0888_ ), .Z(\myreg/_3338_ ) );
BUF_X1 \myreg/_6877_ ( .A(\myreg/_0889_ ), .Z(\myreg/_3339_ ) );
BUF_X1 \myreg/_6878_ ( .A(\myreg/_0890_ ), .Z(\myreg/_3340_ ) );
BUF_X1 \myreg/_6879_ ( .A(\myreg/_0891_ ), .Z(\myreg/_3341_ ) );
BUF_X1 \myreg/_6880_ ( .A(\myreg/_0892_ ), .Z(\myreg/_3342_ ) );
BUF_X1 \myreg/_6881_ ( .A(\myreg/_0893_ ), .Z(\myreg/_3343_ ) );
BUF_X1 \myreg/_6882_ ( .A(\myreg/_0894_ ), .Z(\myreg/_3344_ ) );
BUF_X1 \myreg/_6883_ ( .A(\myreg/_0895_ ), .Z(\myreg/_3345_ ) );
BUF_X1 \myreg/_6884_ ( .A(\myreg/_0896_ ), .Z(\myreg/_3346_ ) );
BUF_X1 \myreg/_6885_ ( .A(\myreg/_0897_ ), .Z(\myreg/_3347_ ) );
BUF_X1 \myreg/_6886_ ( .A(\myreg/_0898_ ), .Z(\myreg/_3348_ ) );
BUF_X1 \myreg/_6887_ ( .A(\myreg/_0899_ ), .Z(\myreg/_3349_ ) );
BUF_X1 \myreg/_6888_ ( .A(\myreg/_0900_ ), .Z(\myreg/_3350_ ) );
BUF_X1 \myreg/_6889_ ( .A(\myreg/_0901_ ), .Z(\myreg/_3351_ ) );
BUF_X1 \myreg/_6890_ ( .A(\myreg/_0902_ ), .Z(\myreg/_3352_ ) );
BUF_X1 \myreg/_6891_ ( .A(\myreg/_0903_ ), .Z(\myreg/_3353_ ) );
BUF_X1 \myreg/_6892_ ( .A(\myreg/_0904_ ), .Z(\myreg/_3354_ ) );
BUF_X1 \myreg/_6893_ ( .A(\myreg/_0905_ ), .Z(\myreg/_3355_ ) );
BUF_X1 \myreg/_6894_ ( .A(\myreg/_0906_ ), .Z(\myreg/_3356_ ) );
BUF_X1 \myreg/_6895_ ( .A(\myreg/_0907_ ), .Z(\myreg/_3357_ ) );
BUF_X1 \myreg/_6896_ ( .A(\myreg/_0908_ ), .Z(\myreg/_3358_ ) );
BUF_X1 \myreg/_6897_ ( .A(\myreg/_0909_ ), .Z(\myreg/_3359_ ) );
BUF_X1 \myreg/_6898_ ( .A(\myreg/_0910_ ), .Z(\myreg/_3360_ ) );
BUF_X1 \myreg/_6899_ ( .A(\myreg/_0911_ ), .Z(\myreg/_3361_ ) );
BUF_X1 \myreg/_6900_ ( .A(\myreg/_0912_ ), .Z(\myreg/_3362_ ) );
BUF_X1 \myreg/_6901_ ( .A(\myreg/_0913_ ), .Z(\myreg/_3363_ ) );
BUF_X1 \myreg/_6902_ ( .A(\myreg/_0914_ ), .Z(\myreg/_3364_ ) );
BUF_X1 \myreg/_6903_ ( .A(\myreg/_0915_ ), .Z(\myreg/_3365_ ) );
BUF_X1 \myreg/_6904_ ( .A(\myreg/_0916_ ), .Z(\myreg/_3366_ ) );
BUF_X1 \myreg/_6905_ ( .A(\myreg/_0917_ ), .Z(\myreg/_3367_ ) );
BUF_X1 \myreg/_6906_ ( .A(\myreg/_0918_ ), .Z(\myreg/_3368_ ) );
BUF_X1 \myreg/_6907_ ( .A(\myreg/_0919_ ), .Z(\myreg/_3369_ ) );
BUF_X1 \myreg/_6908_ ( .A(\myreg/_0920_ ), .Z(\myreg/_3370_ ) );
BUF_X1 \myreg/_6909_ ( .A(\myreg/_0921_ ), .Z(\myreg/_3371_ ) );
BUF_X1 \myreg/_6910_ ( .A(\myreg/_0922_ ), .Z(\myreg/_3372_ ) );
BUF_X1 \myreg/_6911_ ( .A(\myreg/_0923_ ), .Z(\myreg/_3373_ ) );
BUF_X1 \myreg/_6912_ ( .A(\myreg/_0924_ ), .Z(\myreg/_3374_ ) );
BUF_X1 \myreg/_6913_ ( .A(\myreg/_0925_ ), .Z(\myreg/_3375_ ) );
BUF_X1 \myreg/_6914_ ( .A(\myreg/_0926_ ), .Z(\myreg/_3376_ ) );
BUF_X1 \myreg/_6915_ ( .A(\myreg/_0927_ ), .Z(\myreg/_3377_ ) );
BUF_X1 \myreg/_6916_ ( .A(\myreg/_0928_ ), .Z(\myreg/_3378_ ) );
BUF_X1 \myreg/_6917_ ( .A(\myreg/_0929_ ), .Z(\myreg/_3379_ ) );
BUF_X1 \myreg/_6918_ ( .A(\myreg/_0930_ ), .Z(\myreg/_3380_ ) );
BUF_X1 \myreg/_6919_ ( .A(\myreg/_0931_ ), .Z(\myreg/_3381_ ) );
BUF_X1 \myreg/_6920_ ( .A(\myreg/_0932_ ), .Z(\myreg/_3382_ ) );
BUF_X1 \myreg/_6921_ ( .A(\myreg/_0933_ ), .Z(\myreg/_3383_ ) );
BUF_X1 \myreg/_6922_ ( .A(\myreg/_0934_ ), .Z(\myreg/_3384_ ) );
BUF_X1 \myreg/_6923_ ( .A(\myreg/_0935_ ), .Z(\myreg/_3385_ ) );
BUF_X1 \myreg/_6924_ ( .A(\myreg/_0936_ ), .Z(\myreg/_3386_ ) );
BUF_X1 \myreg/_6925_ ( .A(\myreg/_0937_ ), .Z(\myreg/_3387_ ) );
BUF_X1 \myreg/_6926_ ( .A(\myreg/_0938_ ), .Z(\myreg/_3388_ ) );
BUF_X1 \myreg/_6927_ ( .A(\myreg/_0939_ ), .Z(\myreg/_3389_ ) );
BUF_X1 \myreg/_6928_ ( .A(\myreg/_0940_ ), .Z(\myreg/_3390_ ) );
BUF_X1 \myreg/_6929_ ( .A(\myreg/_0941_ ), .Z(\myreg/_3391_ ) );
BUF_X1 \myreg/_6930_ ( .A(\myreg/_0942_ ), .Z(\myreg/_3392_ ) );
BUF_X1 \myreg/_6931_ ( .A(\myreg/_0943_ ), .Z(\myreg/_3393_ ) );
BUF_X1 \myreg/_6932_ ( .A(\myreg/_0944_ ), .Z(\myreg/_3394_ ) );
BUF_X1 \myreg/_6933_ ( .A(\myreg/_0945_ ), .Z(\myreg/_3395_ ) );
BUF_X1 \myreg/_6934_ ( .A(\myreg/_0946_ ), .Z(\myreg/_3396_ ) );
BUF_X1 \myreg/_6935_ ( .A(\myreg/_0947_ ), .Z(\myreg/_3397_ ) );
BUF_X1 \myreg/_6936_ ( .A(\myreg/_0948_ ), .Z(\myreg/_3398_ ) );
BUF_X1 \myreg/_6937_ ( .A(\myreg/_0949_ ), .Z(\myreg/_3399_ ) );
BUF_X1 \myreg/_6938_ ( .A(\myreg/_0950_ ), .Z(\myreg/_3400_ ) );
BUF_X1 \myreg/_6939_ ( .A(\myreg/_0951_ ), .Z(\myreg/_3401_ ) );
BUF_X1 \myreg/_6940_ ( .A(\myreg/_0952_ ), .Z(\myreg/_3402_ ) );
BUF_X1 \myreg/_6941_ ( .A(\myreg/_0953_ ), .Z(\myreg/_3403_ ) );
BUF_X1 \myreg/_6942_ ( .A(\myreg/_0954_ ), .Z(\myreg/_3404_ ) );
BUF_X1 \myreg/_6943_ ( .A(\myreg/_0955_ ), .Z(\myreg/_3405_ ) );
BUF_X1 \myreg/_6944_ ( .A(\myreg/_0956_ ), .Z(\myreg/_3406_ ) );
BUF_X1 \myreg/_6945_ ( .A(\myreg/_0957_ ), .Z(\myreg/_3407_ ) );
BUF_X1 \myreg/_6946_ ( .A(\myreg/_0958_ ), .Z(\myreg/_3408_ ) );
BUF_X1 \myreg/_6947_ ( .A(\myreg/_0959_ ), .Z(\myreg/_3409_ ) );
BUF_X1 \myreg/_6948_ ( .A(\myreg/_0960_ ), .Z(\myreg/_3410_ ) );
BUF_X1 \myreg/_6949_ ( .A(\myreg/_0961_ ), .Z(\myreg/_3411_ ) );
BUF_X1 \myreg/_6950_ ( .A(\myreg/_0962_ ), .Z(\myreg/_3412_ ) );
BUF_X1 \myreg/_6951_ ( .A(\myreg/_0963_ ), .Z(\myreg/_3413_ ) );
BUF_X1 \myreg/_6952_ ( .A(\myreg/_0964_ ), .Z(\myreg/_3414_ ) );
BUF_X1 \myreg/_6953_ ( .A(\myreg/_0965_ ), .Z(\myreg/_3415_ ) );
BUF_X1 \myreg/_6954_ ( .A(\myreg/_0966_ ), .Z(\myreg/_3416_ ) );
BUF_X1 \myreg/_6955_ ( .A(\myreg/_0967_ ), .Z(\myreg/_3417_ ) );
BUF_X1 \myreg/_6956_ ( .A(\myreg/_0968_ ), .Z(\myreg/_3418_ ) );
BUF_X1 \myreg/_6957_ ( .A(\myreg/_0969_ ), .Z(\myreg/_3419_ ) );
BUF_X1 \myreg/_6958_ ( .A(\myreg/_0970_ ), .Z(\myreg/_3420_ ) );
BUF_X1 \myreg/_6959_ ( .A(\myreg/_0971_ ), .Z(\myreg/_3421_ ) );
BUF_X1 \myreg/_6960_ ( .A(\myreg/_0972_ ), .Z(\myreg/_3422_ ) );
BUF_X1 \myreg/_6961_ ( .A(\myreg/_0973_ ), .Z(\myreg/_3423_ ) );
BUF_X1 \myreg/_6962_ ( .A(\myreg/_0974_ ), .Z(\myreg/_3424_ ) );
BUF_X1 \myreg/_6963_ ( .A(\myreg/_0975_ ), .Z(\myreg/_3425_ ) );
BUF_X1 \myreg/_6964_ ( .A(\myreg/_0976_ ), .Z(\myreg/_3426_ ) );
BUF_X1 \myreg/_6965_ ( .A(\myreg/_0977_ ), .Z(\myreg/_3427_ ) );
BUF_X1 \myreg/_6966_ ( .A(\myreg/_0978_ ), .Z(\myreg/_3428_ ) );
BUF_X1 \myreg/_6967_ ( .A(\myreg/_0979_ ), .Z(\myreg/_3429_ ) );
BUF_X1 \myreg/_6968_ ( .A(\myreg/_0980_ ), .Z(\myreg/_3430_ ) );
BUF_X1 \myreg/_6969_ ( .A(\myreg/_0981_ ), .Z(\myreg/_3431_ ) );
BUF_X1 \myreg/_6970_ ( .A(\myreg/_0982_ ), .Z(\myreg/_3432_ ) );
BUF_X1 \myreg/_6971_ ( .A(\myreg/_0983_ ), .Z(\myreg/_3433_ ) );
BUF_X1 \myreg/_6972_ ( .A(\myreg/_0984_ ), .Z(\myreg/_3434_ ) );
BUF_X1 \myreg/_6973_ ( .A(\myreg/_0985_ ), .Z(\myreg/_3435_ ) );
BUF_X1 \myreg/_6974_ ( .A(\myreg/_0986_ ), .Z(\myreg/_3436_ ) );
BUF_X1 \myreg/_6975_ ( .A(\myreg/_0987_ ), .Z(\myreg/_3437_ ) );
BUF_X1 \myreg/_6976_ ( .A(\myreg/_0988_ ), .Z(\myreg/_3438_ ) );
BUF_X1 \myreg/_6977_ ( .A(\myreg/_0989_ ), .Z(\myreg/_3439_ ) );
BUF_X1 \myreg/_6978_ ( .A(\myreg/_0990_ ), .Z(\myreg/_3440_ ) );
BUF_X1 \myreg/_6979_ ( .A(\myreg/_0991_ ), .Z(\myreg/_3441_ ) );
BUF_X1 \myreg/_6980_ ( .A(\myreg/_0992_ ), .Z(\myreg/_3442_ ) );
BUF_X1 \myreg/_6981_ ( .A(\myreg/_0993_ ), .Z(\myreg/_3443_ ) );
BUF_X1 \myreg/_6982_ ( .A(\myreg/_0994_ ), .Z(\myreg/_3444_ ) );
BUF_X1 \myreg/_6983_ ( .A(\myreg/_0995_ ), .Z(\myreg/_3445_ ) );
BUF_X1 \myreg/_6984_ ( .A(\myreg/_0996_ ), .Z(\myreg/_3446_ ) );
BUF_X1 \myreg/_6985_ ( .A(\myreg/_0997_ ), .Z(\myreg/_3447_ ) );
BUF_X1 \myreg/_6986_ ( .A(\myreg/_0998_ ), .Z(\myreg/_3448_ ) );
BUF_X1 \myreg/_6987_ ( .A(\myreg/_0999_ ), .Z(\myreg/_3449_ ) );
BUF_X1 \myreg/_6988_ ( .A(\myreg/_1000_ ), .Z(\myreg/_3450_ ) );
BUF_X1 \myreg/_6989_ ( .A(\myreg/_1001_ ), .Z(\myreg/_3451_ ) );
BUF_X1 \myreg/_6990_ ( .A(\myreg/_1002_ ), .Z(\myreg/_3452_ ) );
BUF_X1 \myreg/_6991_ ( .A(\myreg/_1003_ ), .Z(\myreg/_3453_ ) );
BUF_X1 \myreg/_6992_ ( .A(\myreg/_1004_ ), .Z(\myreg/_3454_ ) );
BUF_X1 \myreg/_6993_ ( .A(\myreg/_1005_ ), .Z(\myreg/_3455_ ) );
BUF_X1 \myreg/_6994_ ( .A(\myreg/_1006_ ), .Z(\myreg/_3456_ ) );
BUF_X1 \myreg/_6995_ ( .A(\myreg/_1007_ ), .Z(\myreg/_3457_ ) );
BUF_X1 \myreg/_6996_ ( .A(\myreg/_1008_ ), .Z(\myreg/_3458_ ) );
BUF_X1 \myreg/_6997_ ( .A(\myreg/_1009_ ), .Z(\myreg/_3459_ ) );
BUF_X1 \myreg/_6998_ ( .A(\myreg/_1010_ ), .Z(\myreg/_3460_ ) );
BUF_X1 \myreg/_6999_ ( .A(\myreg/_1011_ ), .Z(\myreg/_3461_ ) );
BUF_X1 \myreg/_7000_ ( .A(\myreg/_1012_ ), .Z(\myreg/_3462_ ) );
BUF_X1 \myreg/_7001_ ( .A(\myreg/_1013_ ), .Z(\myreg/_3463_ ) );
BUF_X1 \myreg/_7002_ ( .A(\myreg/_1014_ ), .Z(\myreg/_3464_ ) );
BUF_X1 \myreg/_7003_ ( .A(\myreg/_1015_ ), .Z(\myreg/_3465_ ) );
BUF_X1 \myreg/_7004_ ( .A(\myreg/_1016_ ), .Z(\myreg/_3466_ ) );
BUF_X1 \myreg/_7005_ ( .A(\myreg/_1017_ ), .Z(\myreg/_3467_ ) );
BUF_X1 \myreg/_7006_ ( .A(\myreg/_1018_ ), .Z(\myreg/_3468_ ) );
BUF_X1 \myreg/_7007_ ( .A(\myreg/_1019_ ), .Z(\myreg/_3469_ ) );
BUF_X1 \myreg/_7008_ ( .A(\myreg/_1020_ ), .Z(\myreg/_3470_ ) );
BUF_X1 \myreg/_7009_ ( .A(\myreg/_1021_ ), .Z(\myreg/_3471_ ) );
BUF_X1 \myreg/_7010_ ( .A(\myreg/_1022_ ), .Z(\myreg/_3472_ ) );
BUF_X1 \myreg/_7011_ ( .A(\myreg/_1023_ ), .Z(\myreg/_3473_ ) );
INV_X1 \mysc/_28_ ( .A(\mysc/_18_ ), .ZN(\mysc/_10_ ) );
AND3_X1 \mysc/_29_ ( .A1(\mysc/_10_ ), .A2(\mysc/_17_ ), .A3(\mysc/_22_ ), .ZN(\mysc/_05_ ) );
INV_X1 \mysc/_30_ ( .A(\mysc/_20_ ), .ZN(\mysc/_11_ ) );
XOR2_X2 \mysc/_31_ ( .A(\mysc/_03_ ), .B(\mysc/_04_ ), .Z(\mysc/_12_ ) );
AOI21_X1 \mysc/_32_ ( .A(\mysc/_11_ ), .B1(\mysc/_12_ ), .B2(\mysc/_19_ ), .ZN(\mysc/_13_ ) );
OR3_X1 \mysc/_33_ ( .A1(\mysc/_13_ ), .A2(\mysc/_18_ ), .A3(\mysc/_21_ ), .ZN(\mysc/_06_ ) );
NAND4_X1 \mysc/_34_ ( .A1(\mysc/_12_ ), .A2(\mysc/_10_ ), .A3(\mysc/_19_ ), .A4(\mysc/_20_ ), .ZN(\mysc/_14_ ) );
NAND2_X1 \mysc/_35_ ( .A1(\mysc/_10_ ), .A2(\mysc/_22_ ), .ZN(\mysc/_15_ ) );
OAI21_X1 \mysc/_36_ ( .A(\mysc/_14_ ), .B1(\mysc/_17_ ), .B2(\mysc/_15_ ), .ZN(\mysc/_07_ ) );
AND3_X1 \mysc/_37_ ( .A1(\mysc/_10_ ), .A2(\mysc/_22_ ), .A3(\mysc/_09_ ), .ZN(\mysc/_16_ ) );
OR2_X1 \mysc/_38_ ( .A1(\mysc/_05_ ), .A2(\mysc/_16_ ), .ZN(\mysc/_08_ ) );
DFF_X1 \mysc/_39_ ( .D(\mysc/_01_ ), .CK(clock ), .Q(\mysc/state [0] ), .QN(\mysc/_25_ ) );
DFF_X1 \mysc/_40_ ( .D(\mysc/_00_ ), .CK(clock ), .Q(\mysc/state [1] ), .QN(\mysc/_26_ ) );
DFF_X1 \mysc/_41_ ( .D(\mysc/_02_ ), .CK(clock ), .Q(\mysc/state [2] ), .QN(\mysc/_24_ ) );
DFF_X1 \mysc/_42_ ( .D(\mysc/_27_ ), .CK(clock ), .Q(loaduse_clear ), .QN(\mysc/_23_ ) );
BUF_X1 \mysc/_43_ ( .A(reset ), .Z(\mysc/_18_ ) );
BUF_X1 \mysc/_44_ ( .A(previous_load_done ), .Z(\mysc/_17_ ) );
BUF_X1 \mysc/_45_ ( .A(\mysc/state [2] ), .Z(\mysc/_22_ ) );
BUF_X1 \mysc/_46_ ( .A(\mysc/_05_ ), .Z(\mysc/_00_ ) );
BUF_X1 \mysc/_47_ ( .A(\mysc/state [1] ), .Z(\mysc/_21_ ) );
BUF_X1 \mysc/_48_ ( .A(\ID_EX_pc [2] ), .Z(\mysc/_03_ ) );
BUF_X1 \mysc/_49_ ( .A(LS_WB_pc ), .Z(\mysc/_04_ ) );
BUF_X1 \mysc/_50_ ( .A(stall_quest_loaduse ), .Z(\mysc/_19_ ) );
BUF_X1 \mysc/_51_ ( .A(\mysc/state [0] ), .Z(\mysc/_20_ ) );
BUF_X1 \mysc/_52_ ( .A(\mysc/_06_ ), .Z(\mysc/_01_ ) );
BUF_X1 \mysc/_53_ ( .A(\mysc/_07_ ), .Z(\mysc/_02_ ) );
BUF_X1 \mysc/_54_ ( .A(loaduse_clear ), .Z(\mysc/_09_ ) );
BUF_X1 \mysc/_55_ ( .A(\mysc/_08_ ), .Z(\mysc/_27_ ) );
BUF_X8 fanout_buf_1 ( .A(_06_ ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(\myclint/_0000_ ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\myclint/_0329_ ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\mycsreg/_0674_ ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\myexu/_2426_ ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\myexu/_2426_ ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\myexu/_2523_ ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\myexu/_2527_ ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\myexu/myalu/_1360_ ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\myexu/myalu/_1360_ ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\myexu/myalu/_1371_ ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\myexu/myalu/_1371_ ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\myexu/myalu/_1382_ ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\myexu/myalu/_1382_ ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\myexu/myalu/_1385_ ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\myexu/myalu/_1385_ ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myexu/myalu/_1386_ ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myifu/_0930_ ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myifu/_0944_ ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myifu/myicache/_0688_ ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myifu/myicache/_1063_ ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myifu/myicache/_1063_ ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myifu/myicache/_1063_ ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myifu/myicache/_1063_ ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\mylsu/_0310_ ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\mylsu/_0911_ ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\mylsu/_0916_ ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myminixbar/_0486_ ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myreg/_2340_ ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myreg/_2340_ ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myreg/_2340_ ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myreg/_2340_ ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myreg/_2340_ ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myreg/_2340_ ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myreg/_2340_ ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myreg/_2340_ ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myreg/_2340_ ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myreg/_2341_ ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myreg/_2341_ ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myreg/_2341_ ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myreg/_2341_ ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myreg/_2341_ ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myreg/_2341_ ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\myreg/_2342_ ), .Z(fanout_net_44 ) );
BUF_X8 fanout_buf_45 ( .A(\myreg/_2344_ ), .Z(fanout_net_45 ) );
BUF_X8 fanout_buf_46 ( .A(\myreg/_2344_ ), .Z(fanout_net_46 ) );
BUF_X8 fanout_buf_47 ( .A(\myreg/_2344_ ), .Z(fanout_net_47 ) );
BUF_X8 fanout_buf_48 ( .A(\myreg/_2344_ ), .Z(fanout_net_48 ) );
BUF_X8 fanout_buf_49 ( .A(\myreg/_2344_ ), .Z(fanout_net_49 ) );
BUF_X8 fanout_buf_50 ( .A(\myreg/_2344_ ), .Z(fanout_net_50 ) );
BUF_X8 fanout_buf_51 ( .A(\myreg/_2344_ ), .Z(fanout_net_51 ) );
BUF_X8 fanout_buf_52 ( .A(\myreg/_2344_ ), .Z(fanout_net_52 ) );
BUF_X8 fanout_buf_53 ( .A(\myreg/_2344_ ), .Z(fanout_net_53 ) );
BUF_X8 fanout_buf_54 ( .A(fanout_net_59 ), .Z(fanout_net_54 ) );
BUF_X8 fanout_buf_55 ( .A(fanout_net_59 ), .Z(fanout_net_55 ) );
BUF_X8 fanout_buf_56 ( .A(\myreg/_2345_ ), .Z(fanout_net_56 ) );
BUF_X8 fanout_buf_57 ( .A(\myreg/_2345_ ), .Z(fanout_net_57 ) );
BUF_X8 fanout_buf_58 ( .A(\myreg/_2345_ ), .Z(fanout_net_58 ) );
BUF_X8 fanout_buf_59 ( .A(\myreg/_2345_ ), .Z(fanout_net_59 ) );
BUF_X8 fanout_buf_60 ( .A(\myreg/_2346_ ), .Z(fanout_net_60 ) );
BUF_X8 fanout_buf_61 ( .A(\myreg/_2412_ ), .Z(fanout_net_61 ) );

endmodule
